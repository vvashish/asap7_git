# BSD 3-Clause License
# 
# Copyright 2021 Lawrence T. Clark, Vinay Vashishtha, or Arizona State
# University
# 
# Redistribution and use in source and binary forms, with or without
# modification, are permitted provided that the following conditions are met:
# 
# 1. Redistributions of source code must retain the above copyright notice,
# this list of conditions and the following disclaimer.
# 
# 2. Redistributions in binary form must reproduce the above copyright
# notice, this list of conditions and the following disclaimer in the
# documentation and/or other materials provided with the distribution.
# 
# 3. Neither the name of the copyright holder nor the names of its
# contributors may be used to endorse or promote products derived from this
# software without specific prior written permission.
# 
# THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
# AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
# IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
# ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE
# LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
# CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
# SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
# INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
# CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
# ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
# POSSIBILITY OF SUCH DAMAGE.

VERSION 5.8 ;
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 


SITE asap7sc6t 
 CLASS CORE ; 
 SIZE 0.216 BY 0.864 ; 
 SYMMETRY Y ; 
END asap7sc6t 


MACRO A2O1A1Ixp33_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN A2O1A1Ixp33_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.464 0.224 0.612 ; 
        RECT 0.072 0.108 0.144 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.4 0.396 0.568 0.468 ; 
        RECT 0.324 0.464 0.472 0.612 ; 
        RECT 0.4 0.252 0.472 0.612 ; 
        RECT 0.324 0.252 0.472 0.324 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.616 0.54 0.78 0.612 ; 
        RECT 0.708 0.252 0.78 0.612 ; 
        RECT 0.616 0.252 0.78 0.324 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.88 0.54 1.068 0.612 ; 
        RECT 0.996 0.32 1.068 0.612 ; 
        RECT 0.86 0.252 1.008 0.4 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.828 0.684 1.26 0.756 ; 
        RECT 1.188 0.108 1.26 0.756 ; 
        RECT 1.044 0.108 1.26 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.396 0.108 0.9 0.18 ; 
      RECT 0.16 0.684 0.684 0.756 ; 
  END 
END A2O1A1Ixp33_ASAP7_6t_SL 


MACRO A2O1A1Ixp5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN A2O1A1Ixp5_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.54 1.008 0.612 ; 
        RECT 0.936 0.424 1.008 0.612 ; 
        RECT 0.072 0.684 0.308 0.756 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.268 0.396 0.704 0.468 ; 
        RECT 0.268 0.252 0.488 0.324 ; 
        RECT 0.268 0.252 0.34 0.468 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.224 0.252 1.372 0.324 ; 
        RECT 1.152 0.396 1.296 0.468 ; 
        RECT 1.224 0.252 1.296 0.468 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.364 0.54 1.512 0.612 ; 
        RECT 1.44 0.396 1.512 0.612 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.26 0.684 1.656 0.756 ; 
        RECT 1.584 0.108 1.656 0.756 ; 
        RECT 1.476 0.108 1.656 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.612 0.252 1.096 0.324 ; 
      RECT 1.024 0.108 1.096 0.324 ; 
      RECT 1.024 0.108 1.352 0.18 ; 
      RECT 0.592 0.684 1.136 0.756 ; 
      RECT 0.376 0.108 0.9 0.18 ; 
  END 
END A2O1A1Ixp5_ASAP7_6t_SL 


MACRO A2O1A1O1Ixp33_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN A2O1A1O1Ixp33_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.54 0.22 0.612 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.42 0.396 0.576 0.468 ; 
        RECT 0.344 0.536 0.492 0.608 ; 
        RECT 0.42 0.252 0.492 0.608 ; 
        RECT 0.344 0.252 0.492 0.324 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.54 0.872 0.612 ; 
        RECT 0.72 0.252 0.872 0.324 ; 
        RECT 0.72 0.252 0.792 0.612 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.148 0.54 1.3 0.612 ; 
        RECT 1.148 0.252 1.3 0.324 ; 
        RECT 1.148 0.252 1.22 0.612 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.504 0.536 1.656 0.608 ; 
        RECT 1.584 0.252 1.656 0.608 ; 
        RECT 1.504 0.252 1.656 0.324 ; 
    END 
  END D 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.692 0.684 1.872 0.756 ; 
        RECT 1.8 0.108 1.872 0.756 ; 
        RECT 1.044 0.108 1.872 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.808 0.684 1.568 0.756 ; 
      RECT 0.376 0.108 0.92 0.18 ; 
      RECT 0.16 0.684 0.684 0.756 ; 
  END 
END A2O1A1O1Ixp33_ASAP7_6t_SL 


MACRO AND2x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND2x2_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.416 0.54 0.564 0.612 ; 
        RECT 0.492 0.252 0.564 0.612 ; 
        RECT 0.416 0.252 0.564 0.324 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.36 0.468 ; 
        RECT 0.072 0.684 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.684 1.224 0.756 ; 
        RECT 1.152 0.108 1.224 0.756 ; 
        RECT 0.808 0.108 1.224 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.396 0.684 0.708 0.756 ; 
      RECT 0.636 0.108 0.708 0.756 ; 
      RECT 0.636 0.396 0.904 0.468 ; 
      RECT 0.396 0.108 0.708 0.18 ; 
  END 
END AND2x2_ASAP7_6t_SL 


MACRO AND2x4_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND2x4_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.108 1.008 0.468 ; 
        RECT 0.072 0.108 1.008 0.18 ; 
        RECT 0.072 0.684 0.272 0.756 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.404 0.572 0.476 ; 
        RECT 0.352 0.54 0.5 0.612 ; 
        RECT 0.428 0.252 0.5 0.612 ; 
        RECT 0.352 0.252 0.5 0.324 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.26 0.684 2.088 0.756 ; 
        RECT 2.016 0.108 2.088 0.756 ; 
        RECT 1.26 0.108 2.088 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.396 0.684 1.132 0.756 ; 
      RECT 1.06 0.532 1.132 0.756 ; 
      RECT 0.756 0.252 0.828 0.756 ; 
      RECT 1.06 0.532 1.224 0.604 ; 
      RECT 1.152 0.34 1.224 0.604 ; 
      RECT 0.612 0.252 0.828 0.324 ; 
  END 
END AND2x4_ASAP7_6t_SL 


MACRO AND2x6_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND2x6_ASAP7_6t_SL 0 0 ; 
  SIZE 2.592 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.928 0.108 1 0.488 ; 
        RECT 0.072 0.108 1 0.18 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.54 0.648 0.612 ; 
        RECT 0.576 0.396 0.648 0.612 ; 
        RECT 0.428 0.396 0.648 0.468 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.592 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.24 0.684 2.52 0.756 ; 
        RECT 2.448 0.108 2.52 0.756 ; 
        RECT 1.24 0.108 2.52 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.684 1.14 0.756 ; 
      RECT 1.068 0.532 1.14 0.756 ; 
      RECT 0.72 0.252 0.792 0.756 ; 
      RECT 1.068 0.532 1.224 0.604 ; 
      RECT 1.152 0.34 1.224 0.604 ; 
      RECT 0.46 0.252 0.792 0.324 ; 
  END 
END AND2x6_ASAP7_6t_SL 


MACRO AND3x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND3x1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.54 0.22 0.612 ; 
        RECT 0.072 0.108 0.144 0.612 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.396 0.576 0.468 ; 
        RECT 0.352 0.54 0.5 0.612 ; 
        RECT 0.428 0.108 0.5 0.612 ; 
        RECT 0.352 0.108 0.5 0.256 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.644 0.54 0.792 0.612 ; 
        RECT 0.72 0.252 0.792 0.612 ; 
        RECT 0.644 0.252 0.792 0.324 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.044 0.684 1.224 0.756 ; 
        RECT 1.152 0.108 1.224 0.756 ; 
        RECT 1.044 0.108 1.224 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.684 0.936 0.756 ; 
      RECT 0.864 0.108 0.936 0.756 ; 
      RECT 0.864 0.396 1.048 0.468 ; 
      RECT 0.612 0.108 0.936 0.18 ; 
  END 
END AND3x1_ASAP7_6t_SL 


MACRO AND3x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND3x2_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.54 0.22 0.612 ; 
        RECT 0.072 0.108 0.144 0.612 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.42 0.396 0.572 0.468 ; 
        RECT 0.344 0.54 0.492 0.612 ; 
        RECT 0.42 0.108 0.492 0.612 ; 
        RECT 0.344 0.108 0.492 0.256 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.632 0.54 0.78 0.612 ; 
        RECT 0.708 0.252 0.78 0.612 ; 
        RECT 0.632 0.252 0.78 0.324 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.684 1.44 0.756 ; 
        RECT 1.368 0.108 1.44 0.756 ; 
        RECT 1.024 0.108 1.44 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.684 0.924 0.756 ; 
      RECT 0.852 0.108 0.924 0.756 ; 
      RECT 0.852 0.396 1.136 0.468 ; 
      RECT 0.592 0.108 0.924 0.18 ; 
  END 
END AND3x2_ASAP7_6t_SL 


MACRO AND3x4_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND3x4_ASAP7_6t_SL 0 0 ; 
  SIZE 3.024 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.752 0.608 2.956 0.756 ; 
        RECT 2.884 0.252 2.956 0.756 ; 
        RECT 2.808 0.252 2.956 0.324 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.568 0.54 2.268 0.612 ; 
        RECT 2.196 0.396 2.268 0.612 ; 
        RECT 1.568 0.396 2.268 0.468 ; 
        RECT 1.568 0.252 1.716 0.468 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.24 0.54 1.44 0.612 ; 
        RECT 1.368 0.324 1.44 0.612 ; 
        RECT 1.068 0.324 1.44 0.396 ; 
        RECT 1.068 0.108 1.14 0.396 ; 
        RECT 0.992 0.108 1.14 0.18 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.024 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.024 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.684 0.848 0.756 ; 
        RECT 0.776 0.572 0.848 0.756 ; 
        RECT 0.776 0.108 0.848 0.276 ; 
        RECT 0.072 0.108 0.848 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.888 0.252 2.412 0.324 ; 
      RECT 2.34 0.108 2.412 0.324 ; 
      RECT 2.34 0.108 2.872 0.18 ; 
      RECT 0.92 0.684 2.584 0.756 ; 
      RECT 2.512 0.252 2.584 0.756 ; 
      RECT 0.92 0.376 0.992 0.756 ; 
      RECT 2.512 0.252 2.68 0.324 ; 
      RECT 1.24 0.108 2.216 0.18 ; 
  END 
END AND3x4_ASAP7_6t_SL 


MACRO AND4x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND4x1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.036 0.608 0.252 0.756 ; 
        RECT 0.036 0.112 0.252 0.26 ; 
        RECT 0.036 0.396 0.208 0.468 ; 
        RECT 0.036 0.112 0.108 0.756 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.324 0.396 0.588 0.468 ; 
        RECT 0.324 0.396 0.472 0.612 ; 
        RECT 0.324 0.108 0.472 0.256 ; 
        RECT 0.324 0.108 0.396 0.612 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.64 0.54 0.792 0.612 ; 
        RECT 0.72 0.252 0.792 0.612 ; 
        RECT 0.544 0.252 0.792 0.324 ; 
        RECT 0.544 0.108 0.692 0.324 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.908 0.54 1.056 0.612 ; 
        RECT 0.908 0.252 1.056 0.324 ; 
        RECT 0.94 0.252 1.012 0.612 ; 
    END 
  END D 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.3 0.684 1.568 0.756 ; 
        RECT 1.3 0.108 1.568 0.18 ; 
        RECT 1.3 0.108 1.372 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.684 1.228 0.756 ; 
      RECT 1.156 0.108 1.228 0.756 ; 
      RECT 0.828 0.108 1.228 0.18 ; 
  END 
END AND4x1_ASAP7_6t_SL 


MACRO AND4x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND4x2_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.456 0.684 1.692 0.756 ; 
        RECT 1.62 0.112 1.692 0.756 ; 
        RECT 1.52 0.396 1.692 0.468 ; 
        RECT 1.544 0.112 1.692 0.184 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.272 0.396 1.42 0.612 ; 
        RECT 1.348 0.108 1.42 0.612 ; 
        RECT 1.244 0.108 1.42 0.256 ; 
        RECT 1.132 0.396 1.42 0.468 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.252 1.172 0.324 ; 
        RECT 1.024 0.108 1.172 0.324 ; 
        RECT 0.936 0.54 1.088 0.612 ; 
        RECT 0.936 0.252 1.008 0.612 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.664 0.54 0.812 0.612 ; 
        RECT 0.664 0.252 0.812 0.324 ; 
        RECT 0.716 0.252 0.788 0.612 ; 
    END 
  END D 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.16 0.684 0.42 0.756 ; 
        RECT 0.348 0.108 0.42 0.756 ; 
        RECT 0.16 0.108 0.42 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.492 0.684 1.332 0.756 ; 
      RECT 0.492 0.108 0.564 0.756 ; 
      RECT 0.492 0.108 0.9 0.18 ; 
  END 
END AND4x2_ASAP7_6t_SL 


MACRO AND5x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND5x1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.068 0.108 0.26 0.18 ; 
        RECT 0.068 0.108 0.14 0.632 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.412 0.54 0.564 0.612 ; 
        RECT 0.492 0.108 0.564 0.612 ; 
        RECT 0.388 0.108 0.564 0.18 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.712 0.108 0.908 0.18 ; 
        RECT 0.636 0.464 0.784 0.612 ; 
        RECT 0.712 0.108 0.784 0.612 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.008 0.108 1.156 0.208 ; 
        RECT 0.924 0.264 1.08 0.336 ; 
        RECT 1.008 0.108 1.08 0.336 ; 
        RECT 0.856 0.464 1.004 0.612 ; 
        RECT 0.924 0.264 0.996 0.612 ; 
    END 
  END D 
  PIN E 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.18 0.288 1.356 0.36 ; 
        RECT 1.18 0.54 1.336 0.612 ; 
        RECT 1.18 0.288 1.252 0.612 ; 
    END 
  END E 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.592 0.108 1.664 0.656 ; 
        RECT 1.456 0.108 1.664 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.212 0.684 1.508 0.756 ; 
      RECT 1.436 0.384 1.508 0.756 ; 
      RECT 0.212 0.364 0.284 0.756 ; 
      RECT 0.212 0.364 0.36 0.436 ; 
      RECT 0.288 0.264 0.36 0.436 ; 
  END 
END AND5x1_ASAP7_6t_SL 


MACRO AND5x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND5x2_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.068 0.54 0.216 0.612 ; 
        RECT 0.144 0.112 0.216 0.612 ; 
        RECT 0.068 0.112 0.216 0.184 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.396 0.576 0.468 ; 
        RECT 0.288 0.54 0.508 0.612 ; 
        RECT 0.288 0.108 0.436 0.18 ; 
        RECT 0.288 0.108 0.36 0.612 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.252 0.792 0.488 ; 
        RECT 0.564 0.108 0.792 0.18 ; 
        RECT 0.564 0.252 0.792 0.324 ; 
        RECT 0.564 0.108 0.636 0.324 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.864 0.54 1.016 0.612 ; 
        RECT 0.944 0.324 1.016 0.612 ; 
        RECT 0.864 0.252 0.984 0.4 ; 
    END 
  END D 
  PIN E 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.128 0.54 1.276 0.612 ; 
        RECT 1.128 0.252 1.276 0.324 ; 
        RECT 1.152 0.252 1.224 0.612 ; 
    END 
  END E 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.524 0.684 1.872 0.756 ; 
        RECT 1.8 0.108 1.872 0.756 ; 
        RECT 1.524 0.108 1.872 0.18 ; 
        RECT 1.524 0.536 1.596 0.756 ; 
        RECT 1.524 0.108 1.596 0.328 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.132 0.684 1.448 0.756 ; 
      RECT 1.376 0.108 1.448 0.756 ; 
      RECT 1.024 0.108 1.448 0.18 ; 
  END 
END AND5x2_ASAP7_6t_SL 


MACRO AO211x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO211x1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.456 0.252 0.612 0.324 ; 
        RECT 0.516 0.252 0.588 0.48 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.064 0.54 0.212 0.612 ; 
        RECT 0.14 0.108 0.212 0.612 ; 
        RECT 0.064 0.108 0.212 0.18 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.684 1.136 0.756 ; 
        RECT 1.016 0.608 1.136 0.756 ; 
        RECT 1.016 0.396 1.088 0.756 ; 
        RECT 0.936 0.396 1.088 0.468 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.712 0.54 0.892 0.612 ; 
        RECT 0.712 0.252 0.864 0.324 ; 
        RECT 0.712 0.252 0.784 0.612 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.24 0.684 1.476 0.756 ; 
        RECT 1.404 0.108 1.476 0.756 ; 
        RECT 1.196 0.108 1.476 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.284 0.54 0.432 0.612 ; 
      RECT 0.284 0.108 0.356 0.612 ; 
      RECT 1.16 0.252 1.232 0.492 ; 
      RECT 1.16 0.396 1.304 0.468 ; 
      RECT 1 0.252 1.232 0.324 ; 
      RECT 1 0.108 1.072 0.324 ; 
      RECT 0.284 0.108 1.072 0.18 ; 
      RECT 0.16 0.684 0.756 0.756 ; 
  END 
END AO211x1_ASAP7_6t_SL 


MACRO AO211x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO211x2_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.456 0.252 0.612 0.324 ; 
        RECT 0.516 0.252 0.588 0.528 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.064 0.54 0.212 0.612 ; 
        RECT 0.14 0.2 0.212 0.612 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.032 0.56 1.24 0.756 ; 
        RECT 1.016 0.396 1.088 0.608 ; 
        RECT 0.936 0.396 1.088 0.468 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.712 0.252 1.06 0.324 ; 
        RECT 0.784 0.684 0.932 0.756 ; 
        RECT 0.784 0.536 0.856 0.756 ; 
        RECT 0.712 0.252 0.784 0.608 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.312 0.684 1.648 0.756 ; 
        RECT 1.576 0.108 1.648 0.756 ; 
        RECT 1.312 0.108 1.648 0.18 ; 
        RECT 1.312 0.592 1.384 0.756 ; 
        RECT 1.312 0.108 1.384 0.276 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.284 0.54 0.432 0.612 ; 
      RECT 0.284 0.108 0.356 0.612 ; 
      RECT 1.164 0.396 1.384 0.468 ; 
      RECT 1.164 0.108 1.236 0.468 ; 
      RECT 0.284 0.108 1.236 0.18 ; 
      RECT 0.14 0.684 0.684 0.756 ; 
  END 
END AO211x2_ASAP7_6t_SL 


MACRO AO21x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21x1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.068 0.108 0.272 0.18 ; 
        RECT 0.068 0.108 0.14 0.484 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.532 0.54 0.68 0.612 ; 
        RECT 0.532 0.252 0.68 0.324 ; 
        RECT 0.532 0.252 0.604 0.612 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.804 0.608 0.952 0.756 ; 
        RECT 0.804 0.252 0.952 0.4 ; 
        RECT 0.804 0.252 0.876 0.756 ; 
        RECT 0.732 0.396 0.876 0.468 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.608 1.26 0.756 ; 
        RECT 1.188 0.192 1.26 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.284 0.54 0.432 0.612 ; 
      RECT 0.284 0.26 0.356 0.612 ; 
      RECT 1.044 0.108 1.116 0.488 ; 
      RECT 0.284 0.26 0.444 0.332 ; 
      RECT 0.372 0.108 0.444 0.332 ; 
      RECT 0.372 0.108 1.116 0.18 ; 
      RECT 0.16 0.684 0.704 0.756 ; 
  END 
END AO21x1_ASAP7_6t_SL 


MACRO AO21x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21x2_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.064 0.54 0.212 0.612 ; 
        RECT 0.14 0.108 0.212 0.612 ; 
        RECT 0.064 0.108 0.212 0.18 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.512 0.252 0.912 0.324 ; 
        RECT 0.512 0.54 0.668 0.612 ; 
        RECT 0.512 0.252 0.584 0.612 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.728 0.396 1.092 0.468 ; 
        RECT 0.828 0.396 0.976 0.756 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.192 0.684 1.448 0.756 ; 
        RECT 1.192 0.252 1.292 0.756 ; 
        RECT 1.076 0.576 1.292 0.648 ; 
        RECT 1.044 0.252 1.292 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.36 0.108 0.432 0.632 ; 
      RECT 1.368 0.108 1.44 0.468 ; 
      RECT 0.36 0.108 1.44 0.18 ; 
      RECT 0.508 0.684 0.728 0.756 ; 
      RECT 0.064 0.684 0.272 0.756 ; 
    LAYER M2 ; 
      RECT 0.16 0.684 0.716 0.756 ; 
    LAYER V1 ; 
      RECT 0.612 0.684 0.684 0.756 ; 
      RECT 0.18 0.684 0.252 0.756 ; 
  END 
END AO21x2_ASAP7_6t_SL 


MACRO AO221x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO221x1_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.344 0.396 0.564 0.468 ; 
        RECT 0.344 0.396 0.492 0.612 ; 
        RECT 0.344 0.108 0.492 0.256 ; 
        RECT 0.344 0.108 0.416 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.54 0.244 0.612 ; 
        RECT 0.072 0.108 0.144 0.612 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.456 0.684 1.604 0.756 ; 
        RECT 1.456 0.252 1.604 0.324 ; 
        RECT 1.456 0.252 1.528 0.756 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.912 0.252 1.06 0.324 ; 
        RECT 0.836 0.464 0.984 0.612 ; 
        RECT 0.912 0.252 0.984 0.612 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.616 0.54 0.764 0.612 ; 
        RECT 0.692 0.252 0.764 0.612 ; 
        RECT 0.612 0.252 0.764 0.324 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.888 0.684 2.064 0.756 ; 
        RECT 1.992 0.108 2.064 0.756 ; 
        RECT 1.888 0.108 2.064 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.084 0.54 1.344 0.612 ; 
      RECT 1.272 0.108 1.344 0.612 ; 
      RECT 1.716 0.396 1.892 0.468 ; 
      RECT 1.716 0.108 1.788 0.468 ; 
      RECT 0.592 0.108 1.788 0.18 ; 
      RECT 0.828 0.684 1.352 0.756 ; 
      RECT 0.16 0.684 0.704 0.756 ; 
  END 
END AO221x1_ASAP7_6t_SL 


MACRO AO221x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO221x2_ASAP7_6t_SL 0 0 ; 
  SIZE 2.376 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.344 0.396 0.576 0.468 ; 
        RECT 0.344 0.396 0.492 0.612 ; 
        RECT 0.344 0.108 0.492 0.256 ; 
        RECT 0.344 0.108 0.416 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.54 0.244 0.612 ; 
        RECT 0.072 0.108 0.144 0.612 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.456 0.684 1.604 0.756 ; 
        RECT 1.456 0.252 1.604 0.324 ; 
        RECT 1.456 0.252 1.528 0.756 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.912 0.252 1.06 0.324 ; 
        RECT 0.836 0.464 0.984 0.612 ; 
        RECT 0.912 0.252 0.984 0.612 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.616 0.54 0.764 0.612 ; 
        RECT 0.692 0.252 0.764 0.612 ; 
        RECT 0.612 0.252 0.764 0.324 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.376 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.888 0.684 2.064 0.756 ; 
        RECT 1.992 0.108 2.064 0.756 ; 
        RECT 1.888 0.108 2.064 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.084 0.54 1.344 0.612 ; 
      RECT 1.272 0.108 1.344 0.612 ; 
      RECT 1.716 0.396 1.892 0.468 ; 
      RECT 1.716 0.108 1.788 0.468 ; 
      RECT 0.592 0.108 1.788 0.18 ; 
      RECT 0.828 0.684 1.352 0.756 ; 
      RECT 0.16 0.684 0.704 0.756 ; 
  END 
END AO221x2_ASAP7_6t_SL 


MACRO AO222x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO222x1_ASAP7_6t_SL 0 0 ; 
  SIZE 2.376 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.096 0.54 0.276 0.612 ; 
        RECT 0.204 0.108 0.276 0.612 ; 
        RECT 0.096 0.108 0.276 0.18 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.496 0.54 0.668 0.612 ; 
        RECT 0.496 0.252 0.668 0.324 ; 
        RECT 0.496 0.252 0.568 0.612 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.132 0.396 1.352 0.468 ; 
        RECT 1.28 0.252 1.352 0.468 ; 
        RECT 1.132 0.252 1.352 0.324 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.708 0.396 1.012 0.468 ; 
        RECT 0.94 0.252 1.012 0.468 ; 
        RECT 0.792 0.252 1.012 0.324 ; 
    END 
  END B2 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.432 0.396 1.656 0.468 ; 
        RECT 1.432 0.252 1.656 0.324 ; 
        RECT 1.432 0.252 1.504 0.468 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.76 0.252 1.92 0.4 ; 
        RECT 1.644 0.54 1.872 0.612 ; 
        RECT 1.8 0.252 1.872 0.612 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.376 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.1 0.684 2.34 0.756 ; 
        RECT 2.192 0.608 2.34 0.756 ; 
        RECT 2.192 0.108 2.34 0.256 ; 
        RECT 2.192 0.108 2.264 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.348 0.108 0.42 0.632 ; 
      RECT 2.02 0.108 2.092 0.488 ; 
      RECT 0.348 0.108 2.092 0.18 ; 
      RECT 1.368 0.684 1.872 0.756 ; 
      RECT 1.368 0.54 1.44 0.756 ; 
      RECT 0.844 0.54 1.44 0.612 ; 
      RECT 1.024 0.684 1.236 0.756 ; 
      RECT 0.592 0.684 0.74 0.756 ; 
      RECT 0.072 0.684 0.272 0.756 ; 
    LAYER M2 ; 
      RECT 0.08 0.684 1.148 0.756 ; 
    LAYER V1 ; 
      RECT 1.044 0.684 1.116 0.756 ; 
      RECT 0.612 0.684 0.684 0.756 ; 
      RECT 0.18 0.684 0.252 0.756 ; 
  END 
END AO222x1_ASAP7_6t_SL 


MACRO AO222x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO222x2_ASAP7_6t_SL 0 0 ; 
  SIZE 2.592 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.208 0.396 0.28 0.56 ; 
        RECT 0.064 0.108 0.272 0.256 ; 
        RECT 0.064 0.396 0.28 0.468 ; 
        RECT 0.064 0.108 0.136 0.468 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.496 0.252 0.668 0.324 ; 
        RECT 0.496 0.54 0.648 0.612 ; 
        RECT 0.496 0.252 0.568 0.612 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.132 0.396 1.352 0.468 ; 
        RECT 1.28 0.252 1.352 0.468 ; 
        RECT 1.132 0.252 1.352 0.324 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.728 0.396 1.012 0.468 ; 
        RECT 0.8 0.26 1.012 0.468 ; 
    END 
  END B2 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.432 0.396 1.656 0.468 ; 
        RECT 1.432 0.252 1.656 0.324 ; 
        RECT 1.432 0.252 1.504 0.468 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.76 0.252 1.928 0.4 ; 
        RECT 1.644 0.54 1.872 0.612 ; 
        RECT 1.8 0.252 1.872 0.612 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.592 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.104 0.684 2.52 0.756 ; 
        RECT 2.448 0.108 2.52 0.756 ; 
        RECT 2.176 0.108 2.52 0.18 ; 
        RECT 2.176 0.108 2.248 0.296 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.352 0.108 0.424 0.68 ; 
      RECT 2.032 0.108 2.104 0.468 ; 
      RECT 0.352 0.108 2.104 0.18 ; 
      RECT 1.368 0.684 1.872 0.756 ; 
      RECT 1.368 0.54 1.44 0.756 ; 
      RECT 0.844 0.54 1.44 0.612 ; 
      RECT 0.072 0.684 0.26 0.756 ; 
      RECT 0.072 0.608 0.144 0.756 ; 
      RECT 1.024 0.684 1.236 0.756 ; 
      RECT 0.592 0.684 0.74 0.756 ; 
    LAYER M2 ; 
      RECT 0.08 0.684 1.148 0.756 ; 
    LAYER V1 ; 
      RECT 1.044 0.684 1.116 0.756 ; 
      RECT 0.612 0.684 0.684 0.756 ; 
      RECT 0.18 0.684 0.252 0.756 ; 
  END 
END AO222x2_ASAP7_6t_SL 


MACRO AO22x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO22x1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.124 0.54 0.272 0.612 ; 
        RECT 0.2 0.108 0.272 0.612 ; 
        RECT 0.124 0.108 0.272 0.18 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.42 0.392 0.564 0.464 ; 
        RECT 0.344 0.464 0.492 0.612 ; 
        RECT 0.42 0.108 0.492 0.612 ; 
        RECT 0.344 0.108 0.492 0.256 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.236 0.684 1.384 0.756 ; 
        RECT 1.236 0.252 1.384 0.324 ; 
        RECT 1.236 0.252 1.308 0.756 ; 
        RECT 1.144 0.396 1.308 0.468 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.62 0.54 0.768 0.612 ; 
        RECT 0.696 0.108 0.768 0.612 ; 
        RECT 0.592 0.108 0.768 0.26 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.672 0.684 1.832 0.756 ; 
        RECT 1.76 0.108 1.832 0.756 ; 
        RECT 1.672 0.108 1.832 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.868 0.54 1.016 0.612 ; 
      RECT 0.94 0.108 1.016 0.612 ; 
      RECT 1.496 0.396 1.66 0.468 ; 
      RECT 1.496 0.108 1.568 0.468 ; 
      RECT 0.868 0.216 1.016 0.288 ; 
      RECT 0.94 0.108 1.568 0.18 ; 
      RECT 0.16 0.684 1.136 0.756 ; 
  END 
END AO22x1_ASAP7_6t_SL 


MACRO AO22x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO22x2_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.124 0.54 0.272 0.612 ; 
        RECT 0.2 0.108 0.272 0.612 ; 
        RECT 0.124 0.108 0.272 0.18 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.42 0.392 0.564 0.464 ; 
        RECT 0.344 0.464 0.492 0.612 ; 
        RECT 0.42 0.108 0.492 0.612 ; 
        RECT 0.344 0.108 0.492 0.256 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.236 0.684 1.384 0.756 ; 
        RECT 1.236 0.252 1.384 0.324 ; 
        RECT 1.236 0.252 1.308 0.756 ; 
        RECT 1.144 0.396 1.308 0.468 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.62 0.54 0.768 0.612 ; 
        RECT 0.696 0.108 0.768 0.612 ; 
        RECT 0.592 0.108 0.768 0.26 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.672 0.684 1.836 0.756 ; 
        RECT 1.764 0.108 1.836 0.756 ; 
        RECT 1.672 0.108 1.836 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.868 0.54 1.016 0.612 ; 
      RECT 0.94 0.108 1.016 0.612 ; 
      RECT 1.496 0.396 1.66 0.468 ; 
      RECT 1.496 0.108 1.568 0.468 ; 
      RECT 0.868 0.216 1.016 0.288 ; 
      RECT 0.94 0.108 1.568 0.18 ; 
      RECT 0.16 0.684 1.136 0.756 ; 
  END 
END AO22x2_ASAP7_6t_SL 


MACRO AO311x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO311x1_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.712 0.252 0.888 0.324 ; 
        RECT 0.712 0.252 0.784 0.488 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.54 0.576 0.612 ; 
        RECT 0.504 0.108 0.576 0.612 ; 
        RECT 0.376 0.108 0.576 0.18 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.372 0.468 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A3 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.868 0.54 1.016 0.612 ; 
        RECT 0.944 0.384 1.016 0.612 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.252 1.224 0.584 ; 
        RECT 1.076 0.252 1.224 0.324 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.888 0.684 2.084 0.756 ; 
        RECT 2.012 0.108 2.084 0.756 ; 
        RECT 1.888 0.108 2.084 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.24 0.684 1.44 0.756 ; 
      RECT 1.368 0.108 1.44 0.756 ; 
      RECT 1.368 0.396 1.884 0.468 ; 
      RECT 0.792 0.108 1.44 0.18 ; 
      RECT 0.376 0.684 0.936 0.756 ; 
  END 
END AO311x1_ASAP7_6t_SL 


MACRO AO311x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO311x2_ASAP7_6t_SL 0 0 ; 
  SIZE 2.376 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.252 0.868 0.324 ; 
        RECT 0.72 0.252 0.792 0.488 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.54 0.576 0.612 ; 
        RECT 0.504 0.108 0.576 0.612 ; 
        RECT 0.376 0.108 0.576 0.18 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.372 0.468 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A3 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.868 0.54 1.016 0.612 ; 
        RECT 0.944 0.376 1.016 0.612 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.16 0.252 1.232 0.584 ; 
        RECT 1.084 0.252 1.232 0.324 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.376 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.888 0.684 2.3 0.756 ; 
        RECT 2.228 0.108 2.3 0.756 ; 
        RECT 1.888 0.108 2.3 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.24 0.684 1.44 0.756 ; 
      RECT 1.368 0.108 1.44 0.756 ; 
      RECT 1.368 0.396 1.892 0.468 ; 
      RECT 0.792 0.108 1.44 0.18 ; 
      RECT 0.376 0.684 0.936 0.756 ; 
  END 
END AO311x2_ASAP7_6t_SL 


MACRO AO31x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO31x1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.46 0.252 0.612 0.4 ; 
        RECT 0.392 0.54 0.564 0.612 ; 
        RECT 0.492 0.252 0.564 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.712 0.252 0.888 0.324 ; 
        RECT 0.696 0.54 0.844 0.612 ; 
        RECT 0.712 0.252 0.784 0.612 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.02 0.608 1.168 0.756 ; 
        RECT 1.02 0.396 1.092 0.756 ; 
        RECT 0.924 0.396 1.092 0.468 ; 
    END 
  END A3 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.068 0.108 0.216 0.18 ; 
        RECT 0.068 0.108 0.14 0.632 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.292 0.684 1.44 0.756 ; 
        RECT 1.368 0.108 1.44 0.756 ; 
        RECT 1.22 0.108 1.44 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.22 0.296 0.292 0.632 ; 
      RECT 1.224 0.252 1.296 0.488 ; 
      RECT 0.22 0.296 0.388 0.368 ; 
      RECT 0.316 0.108 0.388 0.368 ; 
      RECT 1.024 0.252 1.296 0.324 ; 
      RECT 1.024 0.108 1.096 0.324 ; 
      RECT 0.316 0.108 1.096 0.18 ; 
      RECT 0.376 0.684 0.92 0.756 ; 
  END 
END AO31x1_ASAP7_6t_SL 


MACRO AO31x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO31x2_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.46 0.252 0.608 0.4 ; 
        RECT 0.392 0.54 0.564 0.612 ; 
        RECT 0.492 0.252 0.564 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.712 0.252 0.86 0.324 ; 
        RECT 0.664 0.54 0.828 0.612 ; 
        RECT 0.712 0.252 0.784 0.612 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.016 0.608 1.24 0.756 ; 
        RECT 1.016 0.396 1.088 0.756 ; 
        RECT 0.924 0.396 1.088 0.468 ; 
    END 
  END A3 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.068 0.108 0.216 0.18 ; 
        RECT 0.068 0.108 0.14 0.632 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.312 0.684 1.648 0.756 ; 
        RECT 1.576 0.108 1.648 0.756 ; 
        RECT 1.312 0.108 1.648 0.18 ; 
        RECT 1.312 0.592 1.384 0.756 ; 
        RECT 1.312 0.108 1.384 0.276 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.22 0.296 0.292 0.632 ; 
      RECT 1.16 0.396 1.38 0.468 ; 
      RECT 1.16 0.108 1.232 0.468 ; 
      RECT 0.22 0.296 0.388 0.368 ; 
      RECT 0.316 0.108 0.388 0.368 ; 
      RECT 0.316 0.108 1.232 0.18 ; 
      RECT 0.376 0.684 0.9 0.756 ; 
  END 
END AO31x2_ASAP7_6t_SL 


MACRO AO321x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO321x1_ASAP7_6t_SL 0 0 ; 
  SIZE 2.376 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.376 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.104 0.684 2.3 0.756 ; 
        RECT 2.228 0.108 2.3 0.756 ; 
        RECT 2.104 0.108 2.3 0.18 ; 
    END 
  END Y 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.6 0.396 0.912 0.468 ; 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.488 ; 
      LAYER V1 ; 
        RECT 0.72 0.396 0.792 0.468 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.364 0.252 0.696 0.324 ; 
      LAYER M1 ; 
        RECT 0.392 0.54 0.576 0.612 ; 
        RECT 0.504 0.108 0.576 0.612 ; 
        RECT 0.376 0.108 0.576 0.18 ; 
      LAYER V1 ; 
        RECT 0.504 0.252 0.576 0.324 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 1.032 0.252 1.344 0.324 ; 
      LAYER M1 ; 
        RECT 1.152 0.228 1.224 0.468 ; 
      LAYER V1 ; 
        RECT 1.152 0.252 1.224 0.324 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 1.248 0.396 1.56 0.468 ; 
      LAYER M1 ; 
        RECT 1.356 0.396 1.576 0.468 ; 
        RECT 1.356 0.252 1.576 0.324 ; 
        RECT 1.356 0.252 1.428 0.468 ; 
      LAYER V1 ; 
        RECT 1.368 0.396 1.44 0.468 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.816 0.54 1.128 0.612 ; 
      LAYER M1 ; 
        RECT 0.888 0.54 1.084 0.612 ; 
        RECT 0.936 0.28 1.008 0.612 ; 
      LAYER V1 ; 
        RECT 0.936 0.54 1.008 0.612 ; 
    END 
  END C 
  OBS 
    LAYER M1 ; 
      RECT 1.26 0.54 1.784 0.612 ; 
      RECT 1.712 0.108 1.784 0.612 ; 
      RECT 1.712 0.396 2.1 0.468 ; 
      RECT 1.4 0.108 1.784 0.18 ; 
      RECT 1.044 0.684 1.584 0.756 ; 
      RECT 0.792 0.108 0.952 0.18 ; 
      RECT 0.376 0.684 0.92 0.756 ; 
    LAYER M2 ; 
      RECT 0.808 0.108 1.784 0.18 ; 
    LAYER V1 ; 
      RECT 1.692 0.108 1.764 0.18 ; 
      RECT 0.828 0.108 0.9 0.18 ; 
  END 
END AO321x1_ASAP7_6t_SL 


MACRO AO321x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO321x2_ASAP7_6t_SL 0 0 ; 
  SIZE 2.592 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.592 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.488 ; 
      LAYER M2 ; 
        RECT 0.6 0.396 0.912 0.468 ; 
      LAYER V1 ; 
        RECT 0.72 0.396 0.792 0.468 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.54 0.576 0.612 ; 
        RECT 0.504 0.108 0.576 0.612 ; 
        RECT 0.376 0.108 0.576 0.18 ; 
      LAYER M2 ; 
        RECT 0.384 0.252 0.696 0.324 ; 
      LAYER V1 ; 
        RECT 0.504 0.252 0.576 0.324 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
      LAYER M2 ; 
        RECT 0.072 0.54 0.384 0.612 ; 
      LAYER V1 ; 
        RECT 0.072 0.54 0.144 0.612 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.108 0.108 1.268 0.18 ; 
        RECT 1.152 0.108 1.224 0.468 ; 
      LAYER M2 ; 
        RECT 1.032 0.252 1.344 0.324 ; 
      LAYER V1 ; 
        RECT 1.152 0.252 1.224 0.324 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.356 0.396 1.588 0.468 ; 
        RECT 1.356 0.252 1.588 0.324 ; 
        RECT 1.356 0.252 1.428 0.468 ; 
      LAYER M2 ; 
        RECT 1.32 0.396 1.632 0.468 ; 
      LAYER V1 ; 
        RECT 1.44 0.396 1.512 0.468 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.54 1.084 0.612 ; 
        RECT 0.936 0.28 1.008 0.612 ; 
      LAYER M2 ; 
        RECT 0.824 0.54 1.136 0.612 ; 
      LAYER V1 ; 
        RECT 0.944 0.54 1.016 0.612 ; 
    END 
  END C 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.104 0.684 2.516 0.756 ; 
        RECT 2.444 0.108 2.516 0.756 ; 
        RECT 2.104 0.108 2.516 0.18 ; 
      LAYER M2 ; 
        RECT 2.204 0.396 2.516 0.468 ; 
      LAYER V1 ; 
        RECT 2.444 0.396 2.516 0.468 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.26 0.54 1.784 0.612 ; 
      RECT 1.712 0.108 1.784 0.612 ; 
      RECT 1.712 0.396 2.1 0.468 ; 
      RECT 1.424 0.108 1.784 0.18 ; 
      RECT 1.024 0.684 1.584 0.756 ; 
      RECT 0.792 0.108 0.952 0.18 ; 
      RECT 0.376 0.684 0.9 0.756 ; 
    LAYER M2 ; 
      RECT 0.828 0.108 1.764 0.18 ; 
    LAYER V1 ; 
      RECT 1.692 0.108 1.764 0.18 ; 
      RECT 0.828 0.108 0.9 0.18 ; 
  END 
END AO321x2_ASAP7_6t_SL 


MACRO AO322x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO322x1_ASAP7_6t_SL 0 0 ; 
  SIZE 2.592 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.088 0.464 2.236 0.612 ; 
        RECT 2.016 0.396 2.22 0.468 ; 
        RECT 2.148 0.108 2.22 0.612 ; 
        RECT 2.088 0.384 2.22 0.612 ; 
        RECT 2.072 0.108 2.22 0.256 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.108 2 0.256 ; 
        RECT 1.8 0.54 1.948 0.612 ; 
        RECT 1.8 0.108 1.872 0.612 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.436 0.54 1.7 0.612 ; 
        RECT 1.584 0.108 1.656 0.612 ; 
        RECT 1.484 0.108 1.656 0.256 ; 
        RECT 1.456 0.108 1.656 0.244 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.836 0.396 1.068 0.468 ; 
        RECT 0.996 0.252 1.068 0.468 ; 
        RECT 0.832 0.252 1.068 0.324 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.14 0.396 1.444 0.468 ; 
        RECT 1.14 0.252 1.36 0.324 ; 
        RECT 1.14 0.252 1.212 0.468 ; 
    END 
  END B2 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.068 0.108 0.272 0.256 ; 
        RECT 0.036 0.464 0.184 0.612 ; 
        RECT 0.068 0.108 0.14 0.612 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.488 0.396 0.712 0.468 ; 
        RECT 0.488 0.252 0.708 0.324 ; 
        RECT 0.488 0.252 0.56 0.468 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.592 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.452 0.108 2.524 0.716 ; 
        RECT 2.32 0.108 2.524 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 2.104 0.684 2.38 0.756 ; 
      RECT 2.308 0.376 2.38 0.756 ; 
      RECT 0.128 0.684 0.364 0.756 ; 
      RECT 0.288 0.388 0.364 0.756 ; 
      RECT 0.344 0.108 0.416 0.46 ; 
      RECT 0.344 0.108 1.332 0.18 ; 
      RECT 0.436 0.54 0.508 0.704 ; 
      RECT 0.436 0.54 1.312 0.612 ; 
      RECT 1.044 0.684 1.98 0.756 ; 
      RECT 0.772 0.684 0.92 0.756 ; 
    LAYER M2 ; 
      RECT 0.16 0.684 2.216 0.756 ; 
    LAYER V1 ; 
      RECT 2.124 0.684 2.196 0.756 ; 
      RECT 0.828 0.684 0.9 0.756 ; 
      RECT 0.18 0.684 0.252 0.756 ; 
  END 
END AO322x1_ASAP7_6t_SL 


MACRO AO322x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO322x2_ASAP7_6t_SL 0 0 ; 
  SIZE 2.808 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.152 0.108 2.468 0.18 ; 
        RECT 2.152 0.54 2.316 0.612 ; 
        RECT 2.152 0.108 2.224 0.612 ; 
        RECT 1.996 0.396 2.224 0.468 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.54 2.02 0.612 ; 
        RECT 1.8 0.252 2.02 0.324 ; 
        RECT 1.8 0.252 1.872 0.612 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.656 0.108 2.024 0.18 ; 
        RECT 1.656 0.108 1.728 0.376 ; 
        RECT 1.436 0.54 1.7 0.612 ; 
        RECT 1.584 0.268 1.656 0.612 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.856 0.396 1.076 0.468 ; 
        RECT 1.004 0.252 1.076 0.468 ; 
        RECT 0.856 0.252 1.076 0.324 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.148 0.396 1.444 0.468 ; 
        RECT 1.148 0.252 1.368 0.324 ; 
        RECT 1.148 0.252 1.22 0.468 ; 
    END 
  END B2 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.068 0.54 0.216 0.612 ; 
        RECT 0.144 0.108 0.216 0.612 ; 
        RECT 0.068 0.108 0.216 0.324 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.436 0.396 0.724 0.468 ; 
        RECT 0.436 0.252 0.724 0.324 ; 
        RECT 0.436 0.252 0.508 0.468 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.808 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.808 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.324 0.252 2.74 0.324 ; 
        RECT 2.592 0.108 2.74 0.324 ; 
        RECT 2.268 0.684 2.488 0.756 ; 
        RECT 2.416 0.252 2.488 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 2.604 0.684 2.752 0.756 ; 
      RECT 2.68 0.396 2.752 0.756 ; 
      RECT 2.588 0.396 2.752 0.468 ; 
      RECT 0.144 0.684 0.364 0.756 ; 
      RECT 0.292 0.108 0.364 0.756 ; 
      RECT 0.292 0.108 1.548 0.18 ; 
      RECT 0.448 0.54 0.52 0.704 ; 
      RECT 0.448 0.54 1.312 0.612 ; 
      RECT 1.044 0.684 2 0.756 ; 
      RECT 0.664 0.684 0.92 0.756 ; 
    LAYER M2 ; 
      RECT 0.144 0.684 2.728 0.756 ; 
    LAYER V1 ; 
      RECT 2.628 0.684 2.7 0.756 ; 
      RECT 0.828 0.684 0.9 0.756 ; 
      RECT 0.18 0.684 0.252 0.756 ; 
  END 
END AO322x2_ASAP7_6t_SL 


MACRO AO32x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO32x1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.856 0.464 1.004 0.612 ; 
        RECT 0.932 0.108 1.004 0.612 ; 
        RECT 0.856 0.108 1.004 0.256 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.636 0.464 0.784 0.612 ; 
        RECT 0.712 0.108 0.784 0.612 ; 
        RECT 0.612 0.108 0.784 0.18 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
        RECT 0.492 0.252 0.564 0.612 ; 
        RECT 0.396 0.54 0.564 0.612 ; 
        RECT 0.34 0.608 0.488 0.756 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.076 0.464 1.224 0.612 ; 
        RECT 1.152 0.348 1.224 0.612 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.544 0.108 1.692 0.336 ; 
        RECT 1.516 0.54 1.664 0.612 ; 
        RECT 1.516 0.256 1.588 0.612 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.092 0.684 0.24 0.756 ; 
        RECT 0.092 0.164 0.164 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.296 0.108 1.368 0.64 ; 
      RECT 1.204 0.108 1.444 0.18 ; 
      RECT 0.256 0.108 0.328 0.468 ; 
      RECT 0.256 0.108 0.488 0.18 ; 
      RECT 1.452 0.684 1.664 0.756 ; 
      RECT 0.612 0.684 1.148 0.756 ; 
    LAYER M2 ; 
      RECT 0.808 0.684 1.58 0.756 ; 
      RECT 0.376 0.108 1.412 0.18 ; 
    LAYER V1 ; 
      RECT 1.476 0.684 1.548 0.756 ; 
      RECT 1.26 0.108 1.332 0.18 ; 
      RECT 0.828 0.684 0.9 0.756 ; 
      RECT 0.396 0.108 0.468 0.18 ; 
  END 
END AO32x1_ASAP7_6t_SL 


MACRO AO32x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO32x2_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.072 0.464 1.22 0.612 ; 
        RECT 1.148 0.168 1.22 0.612 ; 
        RECT 1.072 0.168 1.22 0.316 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.852 0.464 1 0.612 ; 
        RECT 0.928 0.176 1 0.612 ; 
        RECT 0.852 0.176 1 0.324 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.552 0.54 0.78 0.612 ; 
        RECT 0.708 0.232 0.78 0.612 ; 
        RECT 0.38 0.684 0.696 0.756 ; 
        RECT 0.552 0.54 0.696 0.756 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.292 0.464 1.44 0.612 ; 
        RECT 1.368 0.168 1.44 0.612 ; 
        RECT 1.292 0.168 1.44 0.316 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.656 0.464 1.88 0.612 ; 
        RECT 1.808 0.252 1.88 0.612 ; 
        RECT 1.684 0.252 1.88 0.34 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.252 0.448 0.324 ; 
        RECT 0.072 0.54 0.428 0.612 ; 
        RECT 0.072 0.54 0.22 0.756 ; 
        RECT 0.072 0.108 0.22 0.324 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.512 0.108 1.584 0.64 ; 
      RECT 1.512 0.108 1.784 0.18 ; 
      RECT 0.336 0.396 0.62 0.468 ; 
      RECT 0.548 0.108 0.62 0.468 ; 
      RECT 0.376 0.108 0.624 0.18 ; 
      RECT 1.672 0.684 1.88 0.756 ; 
      RECT 0.828 0.684 1.364 0.756 ; 
    LAYER M2 ; 
      RECT 1.24 0.684 1.796 0.756 ; 
      RECT 0.376 0.108 1.784 0.18 ; 
    LAYER V1 ; 
      RECT 1.692 0.108 1.764 0.18 ; 
      RECT 1.692 0.684 1.764 0.756 ; 
      RECT 1.26 0.684 1.332 0.756 ; 
      RECT 0.396 0.108 0.468 0.18 ; 
  END 
END AO32x2_ASAP7_6t_SL 


MACRO AO331x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO331x1_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.54 1.084 0.612 ; 
        RECT 0.896 0.108 1.044 0.18 ; 
        RECT 0.936 0.108 1.008 0.612 ; 
      LAYER M2 ; 
        RECT 0.82 0.54 1.204 0.612 ; 
      LAYER V1 ; 
        RECT 0.988 0.54 1.06 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.684 0.54 0.832 0.612 ; 
        RECT 0.724 0.108 0.796 0.612 ; 
        RECT 0.648 0.108 0.796 0.18 ; 
      LAYER M2 ; 
        RECT 0.524 0.396 0.988 0.468 ; 
      LAYER V1 ; 
        RECT 0.724 0.396 0.796 0.468 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.416 0.54 0.576 0.612 ; 
        RECT 0.504 0.396 0.576 0.612 ; 
      LAYER M2 ; 
        RECT 0.304 0.54 0.692 0.612 ; 
      LAYER V1 ; 
        RECT 0.468 0.54 0.54 0.612 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.144 0.108 1.292 0.18 ; 
        RECT 1.144 0.108 1.216 0.44 ; 
      LAYER M2 ; 
        RECT 0.956 0.252 1.42 0.324 ; 
      LAYER V1 ; 
        RECT 1.144 0.252 1.216 0.324 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.336 0.396 1.484 0.468 ; 
        RECT 1.372 0.28 1.444 0.468 ; 
      LAYER M2 ; 
        RECT 1.172 0.396 1.648 0.468 ; 
      LAYER V1 ; 
        RECT 1.388 0.396 1.46 0.468 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.252 1.772 0.324 ; 
        RECT 1.584 0.252 1.656 0.44 ; 
      LAYER M2 ; 
        RECT 1.608 0.252 2.044 0.324 ; 
      LAYER V1 ; 
        RECT 1.692 0.252 1.764 0.324 ; 
    END 
  END B3 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.808 0.396 1.98 0.468 ; 
        RECT 1.908 0.28 1.98 0.468 ; 
      LAYER M2 ; 
        RECT 1.784 0.396 2.044 0.468 ; 
      LAYER V1 ; 
        RECT 1.876 0.396 1.948 0.468 ; 
    END 
  END C 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.684 0.272 0.756 ; 
        RECT 0.072 0.108 0.252 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
      LAYER M2 ; 
        RECT 0.156 0.684 0.548 0.756 ; 
      LAYER V1 ; 
        RECT 0.18 0.684 0.252 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.808 0.684 2.124 0.756 ; 
      RECT 2.052 0.108 2.124 0.756 ; 
      RECT 1.456 0.108 2.124 0.18 ; 
      RECT 0.288 0.252 0.36 0.468 ; 
      RECT 0.288 0.252 0.448 0.324 ; 
      RECT 0.376 0.108 0.448 0.324 ; 
      RECT 0.376 0.108 0.524 0.18 ; 
      RECT 1.26 0.54 1.86 0.612 ; 
      RECT 0.552 0.684 1.572 0.756 ; 
    LAYER M2 ; 
      RECT 0.376 0.108 1.784 0.18 ; 
    LAYER V1 ; 
      RECT 1.692 0.108 1.764 0.18 ; 
      RECT 0.396 0.108 0.468 0.18 ; 
  END 
END AO331x1_ASAP7_6t_SL 


MACRO AO331x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO331x2_ASAP7_6t_SL 0 0 ; 
  SIZE 2.376 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.376 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.54 1.308 0.612 ; 
        RECT 1.152 0.212 1.224 0.612 ; 
      LAYER M2 ; 
        RECT 1.052 0.54 1.52 0.612 ; 
      LAYER V1 ; 
        RECT 1.188 0.54 1.26 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.9 0.54 1.048 0.612 ; 
        RECT 0.932 0.212 1.004 0.612 ; 
      LAYER M2 ; 
        RECT 0.824 0.252 1.12 0.324 ; 
      LAYER V1 ; 
        RECT 0.932 0.252 1.004 0.324 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.644 0.54 0.792 0.612 ; 
        RECT 0.72 0.396 0.792 0.612 ; 
      LAYER M2 ; 
        RECT 0.452 0.54 0.896 0.612 ; 
      LAYER V1 ; 
        RECT 0.668 0.54 0.74 0.612 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.344 0.396 1.456 0.468 ; 
        RECT 1.36 0.212 1.432 0.468 ; 
      LAYER M2 ; 
        RECT 1.34 0.396 1.648 0.468 ; 
      LAYER V1 ; 
        RECT 1.368 0.396 1.44 0.468 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.532 0.252 1.7 0.324 ; 
        RECT 1.588 0.252 1.66 0.44 ; 
      LAYER M2 ; 
        RECT 1.532 0.252 1.812 0.324 ; 
      LAYER V1 ; 
        RECT 1.552 0.252 1.624 0.324 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.252 2.136 0.324 ; 
        RECT 1.8 0.252 1.872 0.44 ; 
      LAYER M2 ; 
        RECT 1.936 0.252 2.288 0.324 ; 
      LAYER V1 ; 
        RECT 2.016 0.252 2.088 0.324 ; 
    END 
  END B3 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.996 0.396 2.168 0.468 ; 
      LAYER M2 ; 
        RECT 1.936 0.396 2.288 0.468 ; 
      LAYER V1 ; 
        RECT 2.016 0.396 2.088 0.468 ; 
    END 
  END C 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.684 0.488 0.756 ; 
        RECT 0.072 0.108 0.468 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
      LAYER M2 ; 
        RECT 0.372 0.684 0.764 0.756 ; 
      LAYER V1 ; 
        RECT 0.396 0.684 0.468 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 2.104 0.684 2.34 0.756 ; 
      RECT 2.268 0.108 2.34 0.756 ; 
      RECT 1.672 0.108 2.34 0.18 ; 
      RECT 0.42 0.252 0.492 0.488 ; 
      RECT 0.42 0.252 0.672 0.324 ; 
      RECT 0.592 0.108 0.672 0.324 ; 
      RECT 0.592 0.108 0.74 0.18 ; 
      RECT 1.496 0.54 2 0.612 ; 
      RECT 0.788 0.684 1.788 0.756 ; 
    LAYER M2 ; 
      RECT 0.592 0.108 1.784 0.18 ; 
    LAYER V1 ; 
      RECT 1.692 0.108 1.764 0.18 ; 
      RECT 0.612 0.108 0.684 0.18 ; 
  END 
END AO331x2_ASAP7_6t_SL 


MACRO AO332x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO332x1_ASAP7_6t_SL 0 0 ; 
  SIZE 3.024 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.636 0.388 0.8 0.46 ; 
        RECT 0.636 0.108 0.708 0.632 ; 
        RECT 0.376 0.108 0.708 0.18 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.54 0.564 0.612 ; 
        RECT 0.492 0.252 0.564 0.612 ; 
        RECT 0.272 0.252 0.564 0.324 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.848 0.54 0.996 0.612 ; 
        RECT 0.924 0.108 0.996 0.612 ; 
        RECT 0.808 0.108 0.996 0.18 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.068 0.108 1.352 0.18 ; 
        RECT 1.068 0.396 1.288 0.468 ; 
        RECT 1.068 0.108 1.14 0.468 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.428 0.396 1.648 0.468 ; 
        RECT 1.24 0.252 1.648 0.324 ; 
        RECT 1.428 0.252 1.5 0.468 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.32 0.684 2.528 0.756 ; 
        RECT 2.456 0.252 2.528 0.756 ; 
        RECT 2.368 0.252 2.528 0.324 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.78 0.396 2.12 0.468 ; 
        RECT 2.048 0.252 2.12 0.468 ; 
        RECT 1.78 0.252 2.12 0.324 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.024 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.024 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.752 0.684 2.952 0.756 ; 
        RECT 2.88 0.108 2.952 0.756 ; 
        RECT 2.804 0.108 2.952 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.928 0.54 2.268 0.612 ; 
      RECT 2.196 0.108 2.268 0.612 ; 
      RECT 2.6 0.396 2.78 0.468 ; 
      RECT 2.6 0.108 2.672 0.468 ; 
      RECT 1.476 0.108 2.672 0.18 ; 
      RECT 1.732 0.684 2.196 0.756 ; 
      RECT 1.732 0.54 1.804 0.756 ; 
      RECT 1.1 0.54 1.804 0.612 ; 
      RECT 0.772 0.684 1.568 0.756 ; 
      RECT 0.376 0.684 0.54 0.756 ; 
    LAYER M2 ; 
      RECT 0.396 0.684 0.936 0.756 ; 
    LAYER V1 ; 
      RECT 0.828 0.684 0.9 0.756 ; 
      RECT 0.396 0.684 0.468 0.756 ; 
  END 
END AO332x1_ASAP7_6t_SL 


MACRO AO332x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO332x2_ASAP7_6t_SL 0 0 ; 
  SIZE 3.24 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.636 0.388 0.8 0.46 ; 
        RECT 0.636 0.108 0.708 0.632 ; 
        RECT 0.376 0.108 0.708 0.18 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.54 0.564 0.612 ; 
        RECT 0.492 0.252 0.564 0.612 ; 
        RECT 0.272 0.252 0.564 0.324 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.828 0.54 0.996 0.612 ; 
        RECT 0.924 0.108 0.996 0.612 ; 
        RECT 0.808 0.108 0.996 0.18 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.068 0.108 1.352 0.18 ; 
        RECT 1.068 0.396 1.288 0.468 ; 
        RECT 1.068 0.108 1.14 0.468 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.428 0.396 1.648 0.468 ; 
        RECT 1.24 0.252 1.648 0.324 ; 
        RECT 1.428 0.252 1.5 0.468 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.32 0.684 2.528 0.756 ; 
        RECT 2.456 0.252 2.528 0.756 ; 
        RECT 2.368 0.252 2.528 0.324 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.78 0.396 2.12 0.468 ; 
        RECT 2.048 0.252 2.12 0.468 ; 
        RECT 1.78 0.252 2.12 0.324 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.24 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.24 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.808 0.684 3.168 0.756 ; 
        RECT 3.096 0.108 3.168 0.756 ; 
        RECT 2.804 0.108 3.168 0.18 ; 
        RECT 2.808 0.592 2.88 0.756 ; 
        RECT 2.804 0.108 2.876 0.272 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.928 0.54 2.268 0.612 ; 
      RECT 2.196 0.108 2.268 0.612 ; 
      RECT 2.6 0.396 2.78 0.468 ; 
      RECT 2.6 0.108 2.672 0.468 ; 
      RECT 1.476 0.108 2.672 0.18 ; 
      RECT 1.732 0.684 2.196 0.756 ; 
      RECT 1.732 0.54 1.804 0.756 ; 
      RECT 1.1 0.54 1.804 0.612 ; 
      RECT 0.772 0.684 1.568 0.756 ; 
      RECT 0.376 0.684 0.54 0.756 ; 
    LAYER M2 ; 
      RECT 0.396 0.684 0.936 0.756 ; 
    LAYER V1 ; 
      RECT 0.828 0.684 0.9 0.756 ; 
      RECT 0.396 0.684 0.468 0.756 ; 
  END 
END AO332x2_ASAP7_6t_SL 


MACRO AO333x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO333x1_ASAP7_6t_SL 0 0 ; 
  SIZE 3.456 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.736 0.54 2.884 0.612 ; 
        RECT 2.736 0.252 2.884 0.324 ; 
        RECT 2.736 0.252 2.808 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.516 0.252 2.664 0.612 ; 
        RECT 2.22 0.396 2.664 0.468 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.32 0.108 2.552 0.18 ; 
        RECT 1.864 0.252 2.392 0.324 ; 
        RECT 2.32 0.108 2.392 0.324 ; 
        RECT 1.864 0.396 2.096 0.468 ; 
        RECT 1.864 0.252 1.936 0.468 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.82 0.54 0.996 0.612 ; 
        RECT 0.924 0.108 0.996 0.612 ; 
        RECT 0.808 0.108 0.996 0.18 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.068 0.396 1.288 0.468 ; 
        RECT 1.068 0.108 1.288 0.18 ; 
        RECT 1.068 0.108 1.14 0.636 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.428 0.396 1.668 0.468 ; 
        RECT 1.24 0.252 1.648 0.324 ; 
        RECT 1.428 0.252 1.5 0.468 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.636 0.388 0.8 0.46 ; 
        RECT 0.636 0.108 0.708 0.632 ; 
        RECT 0.376 0.108 0.708 0.18 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.54 0.564 0.612 ; 
        RECT 0.492 0.252 0.564 0.612 ; 
        RECT 0.372 0.252 0.564 0.324 ; 
    END 
  END C2 
  PIN C3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END C3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.456 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.456 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 3.184 0.684 3.384 0.756 ; 
        RECT 3.312 0.108 3.384 0.756 ; 
        RECT 3.184 0.108 3.384 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 2.536 0.684 3.056 0.756 ; 
      RECT 2.984 0.528 3.056 0.756 ; 
      RECT 3.028 0.256 3.1 0.608 ; 
      RECT 2.984 0.108 3.056 0.336 ; 
      RECT 2.752 0.108 3.056 0.18 ; 
      RECT 2.34 0.54 2.412 0.704 ; 
      RECT 1.252 0.54 1.324 0.704 ; 
      RECT 1.252 0.54 2.412 0.612 ; 
      RECT 2.02 0.684 2.216 0.756 ; 
      RECT 1.456 0.108 2.196 0.18 ; 
      RECT 1.452 0.684 1.652 0.756 ; 
      RECT 0.772 0.684 0.956 0.756 ; 
      RECT 0.376 0.684 0.54 0.756 ; 
    LAYER M2 ; 
      RECT 2.084 0.684 2.72 0.756 ; 
      RECT 0.396 0.684 1.62 0.756 ; 
    LAYER V1 ; 
      RECT 2.556 0.684 2.628 0.756 ; 
      RECT 2.124 0.684 2.196 0.756 ; 
      RECT 1.476 0.684 1.548 0.756 ; 
      RECT 0.828 0.684 0.9 0.756 ; 
      RECT 0.396 0.684 0.468 0.756 ; 
  END 
END AO333x1_ASAP7_6t_SL 


MACRO AO333x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO333x2_ASAP7_6t_SL 0 0 ; 
  SIZE 3.672 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.736 0.54 2.884 0.612 ; 
        RECT 2.736 0.252 2.884 0.324 ; 
        RECT 2.736 0.252 2.808 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.516 0.252 2.664 0.612 ; 
        RECT 2.22 0.396 2.664 0.468 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.32 0.108 2.552 0.18 ; 
        RECT 1.864 0.252 2.392 0.324 ; 
        RECT 2.32 0.108 2.392 0.324 ; 
        RECT 1.864 0.396 2.088 0.468 ; 
        RECT 1.864 0.252 1.936 0.468 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.82 0.54 0.996 0.612 ; 
        RECT 0.924 0.108 0.996 0.612 ; 
        RECT 0.808 0.108 0.996 0.18 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.068 0.396 1.288 0.468 ; 
        RECT 1.068 0.108 1.288 0.18 ; 
        RECT 1.068 0.108 1.14 0.636 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.428 0.396 1.648 0.468 ; 
        RECT 1.24 0.252 1.648 0.324 ; 
        RECT 1.428 0.252 1.5 0.468 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.636 0.388 0.8 0.46 ; 
        RECT 0.636 0.108 0.708 0.632 ; 
        RECT 0.376 0.108 0.708 0.18 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.54 0.564 0.612 ; 
        RECT 0.492 0.252 0.564 0.612 ; 
        RECT 0.364 0.252 0.564 0.324 ; 
    END 
  END C2 
  PIN C3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.252 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END C3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.672 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.672 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 3.184 0.684 3.384 0.756 ; 
        RECT 3.312 0.108 3.384 0.756 ; 
        RECT 3.184 0.108 3.384 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 2.536 0.684 3.056 0.756 ; 
      RECT 2.984 0.528 3.056 0.756 ; 
      RECT 3.028 0.256 3.1 0.608 ; 
      RECT 2.984 0.108 3.056 0.336 ; 
      RECT 2.752 0.108 3.056 0.18 ; 
      RECT 2.34 0.54 2.412 0.704 ; 
      RECT 1.252 0.54 1.324 0.704 ; 
      RECT 1.252 0.54 2.412 0.612 ; 
      RECT 2.02 0.684 2.216 0.756 ; 
      RECT 1.456 0.108 2.196 0.18 ; 
      RECT 1.452 0.684 1.652 0.756 ; 
      RECT 0.772 0.684 0.956 0.756 ; 
      RECT 0.376 0.684 0.54 0.756 ; 
    LAYER M2 ; 
      RECT 2.084 0.684 2.72 0.756 ; 
      RECT 0.396 0.684 1.62 0.756 ; 
    LAYER V1 ; 
      RECT 2.556 0.684 2.628 0.756 ; 
      RECT 2.124 0.684 2.196 0.756 ; 
      RECT 1.476 0.684 1.548 0.756 ; 
      RECT 0.828 0.684 0.9 0.756 ; 
      RECT 0.396 0.684 0.468 0.756 ; 
  END 
END AO333x2_ASAP7_6t_SL 


MACRO AO33x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO33x1_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.748 0.54 1.008 0.612 ; 
        RECT 0.936 0.108 1.008 0.612 ; 
        RECT 0.808 0.108 1.008 0.256 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.108 0.54 1.268 0.612 ; 
        RECT 1.108 0.252 1.26 0.324 ; 
        RECT 1.152 0.252 1.224 0.612 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.548 0.396 0.812 0.468 ; 
        RECT 0.548 0.108 0.704 0.18 ; 
        RECT 0.548 0.108 0.62 0.68 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.36 0.108 1.432 0.44 ; 
        RECT 1.12 0.108 1.432 0.18 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.504 0.108 1.832 0.18 ; 
        RECT 1.504 0.396 1.668 0.468 ; 
        RECT 1.504 0.108 1.576 0.468 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.94 0.108 2.096 0.18 ; 
        RECT 1.94 0.396 2.088 0.468 ; 
        RECT 1.94 0.108 2.012 0.468 ; 
    END 
  END B3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.284 0.54 0.448 0.612 ; 
        RECT 0.284 0.22 0.448 0.292 ; 
        RECT 0.284 0.108 0.356 0.612 ; 
        RECT 0.16 0.108 0.356 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.9 0.684 2.092 0.756 ; 
      RECT 1.9 0.54 2.016 0.756 ; 
      RECT 1.412 0.54 2.016 0.612 ; 
      RECT 1.796 0.252 1.868 0.612 ; 
      RECT 1.704 0.252 1.868 0.324 ; 
      RECT 0.072 0.684 0.292 0.756 ; 
      RECT 0.072 0.368 0.144 0.756 ; 
      RECT 0.804 0.684 1.764 0.756 ; 
    LAYER M2 ; 
      RECT 0.1 0.684 2.056 0.756 ; 
    LAYER V1 ; 
      RECT 1.908 0.684 1.98 0.756 ; 
      RECT 0.18 0.684 0.252 0.756 ; 
  END 
END AO33x1_ASAP7_6t_SL 


MACRO AO33x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO33x2_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.748 0.54 1.008 0.612 ; 
        RECT 0.936 0.108 1.008 0.612 ; 
        RECT 0.808 0.108 1.008 0.256 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.108 0.54 1.268 0.612 ; 
        RECT 1.108 0.252 1.26 0.324 ; 
        RECT 1.152 0.252 1.224 0.612 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.548 0.396 0.812 0.468 ; 
        RECT 0.548 0.108 0.704 0.256 ; 
        RECT 0.548 0.108 0.62 0.652 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.36 0.108 1.432 0.44 ; 
        RECT 1.12 0.108 1.432 0.18 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.504 0.108 1.782 0.18 ; 
        RECT 1.504 0.396 1.668 0.468 ; 
        RECT 1.504 0.108 1.576 0.468 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.952 0.108 2.124 0.324 ; 
        RECT 2.024 0.108 2.096 0.468 ; 
    END 
  END B3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.404 0.416 0.476 0.652 ; 
        RECT 0.284 0.22 0.448 0.292 ; 
        RECT 0.284 0.416 0.476 0.488 ; 
        RECT 0.284 0.108 0.356 0.488 ; 
        RECT 0.08 0.108 0.356 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.896 0.684 2.088 0.756 ; 
      RECT 1.896 0.54 1.988 0.756 ; 
      RECT 1.412 0.54 1.988 0.612 ; 
      RECT 1.796 0.252 1.868 0.612 ; 
      RECT 1.704 0.252 1.868 0.324 ; 
      RECT 0.072 0.68 0.272 0.756 ; 
      RECT 0.072 0.368 0.144 0.756 ; 
      RECT 0.804 0.684 1.764 0.756 ; 
    LAYER M2 ; 
      RECT 0.1 0.684 2.052 0.756 ; 
    LAYER V1 ; 
      RECT 1.908 0.684 1.98 0.756 ; 
      RECT 0.18 0.684 0.252 0.756 ; 
  END 
END AO33x2_ASAP7_6t_SL 


MACRO AOI211xp25_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI211xp25_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.18 0.576 0.416 ; 
        RECT 0.424 0.18 0.576 0.252 ; 
      LAYER M2 ; 
        RECT 0.252 0.252 0.604 0.324 ; 
      LAYER V1 ; 
        RECT 0.504 0.252 0.576 0.324 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.28 0.144 0.584 ; 
      LAYER M2 ; 
        RECT 0.072 0.396 0.392 0.468 ; 
      LAYER V1 ; 
        RECT 0.072 0.396 0.144 0.468 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.712 0.252 0.86 0.324 ; 
        RECT 0.712 0.252 0.784 0.488 ; 
      LAYER M2 ; 
        RECT 0.692 0.396 1.1 0.468 ; 
      LAYER V1 ; 
        RECT 0.712 0.396 0.784 0.468 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.868 0.54 1.016 0.612 ; 
        RECT 0.944 0.376 1.016 0.612 ; 
      LAYER M2 ; 
        RECT 0.636 0.54 0.972 0.612 ; 
      LAYER V1 ; 
        RECT 0.88 0.54 0.952 0.612 ; 
    END 
  END C 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.988 0.684 1.224 0.756 ; 
        RECT 1.152 0.108 1.224 0.756 ; 
        RECT 0.72 0.108 1.224 0.18 ; 
        RECT 0.252 0.54 0.468 0.612 ; 
        RECT 0.252 0.108 0.324 0.612 ; 
        RECT 0.16 0.108 0.324 0.18 ; 
      LAYER M2 ; 
        RECT 0.16 0.108 1.116 0.18 ; 
      LAYER V1 ; 
        RECT 0.18 0.108 0.252 0.18 ; 
        RECT 1.044 0.108 1.116 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.684 0.704 0.756 ; 
  END 
END AOI211xp25_ASAP7_6t_SL 


MACRO AOI211xp5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI211xp5_ASAP7_6t_SL 0 0 ; 
  SIZE 2.592 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.472 0.468 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.592 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.708 0.396 0.98 0.468 ; 
      LAYER M1 ; 
        RECT 0.636 0.396 0.952 0.468 ; 
        RECT 0.636 0.54 0.936 0.612 ; 
        RECT 0.636 0.108 0.936 0.18 ; 
        RECT 0.636 0.108 0.708 0.612 ; 
      LAYER V1 ; 
        RECT 0.808 0.396 0.88 0.468 ; 
    END 
  END A1 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 1.156 0.252 1.428 0.324 ; 
      LAYER M1 ; 
        RECT 1.256 0.396 1.476 0.468 ; 
        RECT 1.256 0.108 1.476 0.18 ; 
        RECT 1.256 0.108 1.328 0.468 ; 
      LAYER V1 ; 
        RECT 1.256 0.252 1.328 0.324 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 1.98 0.396 2.252 0.468 ; 
      LAYER M1 ; 
        RECT 2.048 0.396 2.268 0.468 ; 
        RECT 2.196 0.252 2.268 0.468 ; 
        RECT 2.048 0.252 2.268 0.324 ; 
      LAYER V1 ; 
        RECT 2.08 0.396 2.152 0.468 ; 
    END 
  END C 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.376 0.108 2.432 0.18 ; 
      LAYER M1 ; 
        RECT 2.076 0.54 2.548 0.612 ; 
        RECT 2.476 0.108 2.548 0.612 ; 
        RECT 2.332 0.108 2.548 0.18 ; 
        RECT 1.812 0.108 2 0.18 ; 
        RECT 0.376 0.108 0.524 0.18 ; 
      LAYER V1 ; 
        RECT 0.396 0.108 0.468 0.18 ; 
        RECT 1.908 0.108 1.98 0.18 ; 
        RECT 2.34 0.108 2.412 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.684 1.224 0.756 ; 
      RECT 1.152 0.54 1.224 0.756 ; 
      RECT 1.152 0.54 1.796 0.612 ; 
      RECT 1.444 0.684 2.432 0.756 ; 
  END 
END AOI211xp5_ASAP7_6t_SL 


MACRO AOI21x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21x1_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.632 0.396 1.332 0.468 ; 
        RECT 0.556 0.54 0.704 0.612 ; 
        RECT 0.632 0.252 0.704 0.612 ; 
        RECT 0.556 0.252 0.704 0.324 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.392 0.308 0.464 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.456 0.396 1.844 0.468 ; 
        RECT 1.772 0.252 1.844 0.468 ; 
        RECT 1.58 0.252 1.844 0.324 ; 
        RECT 1.22 0.54 1.528 0.612 ; 
        RECT 1.456 0.396 1.528 0.612 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.672 0.54 2.056 0.612 ; 
        RECT 1.984 0.108 2.056 0.612 ; 
        RECT 1.024 0.108 2.056 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.828 0.252 1.352 0.324 ; 
      RECT 0.828 0.108 0.9 0.324 ; 
      RECT 0.376 0.108 0.9 0.18 ; 
      RECT 0.376 0.684 2 0.756 ; 
  END 
END AOI21x1_ASAP7_6t_SL 


MACRO AOI21xp25_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21xp25_ASAP7_6t_SL 0 0 ; 
  SIZE 1.08 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.344 0.392 0.584 0.464 ; 
        RECT 0.344 0.108 0.492 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.112 0.464 0.272 0.612 ; 
        RECT 0.112 0.108 0.272 0.288 ; 
        RECT 0.112 0.108 0.184 0.612 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.54 0.868 0.612 ; 
        RECT 0.72 0.252 0.868 0.324 ; 
        RECT 0.72 0.252 0.792 0.612 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.08 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.08 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.684 1.044 0.756 ; 
        RECT 0.972 0.108 1.044 0.756 ; 
        RECT 0.592 0.108 1.044 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.684 0.684 0.756 ; 
  END 
END AOI21xp25_ASAP7_6t_SL 


MACRO AOI21xp5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21xp5_ASAP7_6t_SL 0 0 ; 
  SIZE 1.08 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.344 0.392 0.584 0.464 ; 
        RECT 0.344 0.108 0.492 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.112 0.464 0.272 0.612 ; 
        RECT 0.112 0.108 0.272 0.272 ; 
        RECT 0.112 0.108 0.184 0.612 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.54 0.868 0.612 ; 
        RECT 0.72 0.252 0.868 0.324 ; 
        RECT 0.72 0.252 0.792 0.612 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.08 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.08 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.684 1.044 0.756 ; 
        RECT 0.972 0.108 1.044 0.756 ; 
        RECT 0.592 0.108 1.044 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.684 0.684 0.756 ; 
  END 
END AOI21xp5_ASAP7_6t_SL 


MACRO AOI221xp25_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI221xp25_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.952 0.54 1.172 0.612 ; 
        RECT 1.1 0.108 1.172 0.612 ; 
        RECT 0.936 0.396 1.172 0.468 ; 
        RECT 1.024 0.108 1.172 0.18 ; 
      LAYER M2 ; 
        RECT 0.868 0.54 1.236 0.612 ; 
      LAYER V1 ; 
        RECT 1.008 0.54 1.08 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.244 0.464 1.44 0.612 ; 
        RECT 1.368 0.112 1.44 0.612 ; 
        RECT 1.244 0.112 1.44 0.26 ; 
      LAYER M2 ; 
        RECT 1.184 0.396 1.44 0.468 ; 
      LAYER V1 ; 
        RECT 1.368 0.396 1.44 0.468 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.232 0.144 0.604 ; 
      LAYER M2 ; 
        RECT 0.072 0.396 0.328 0.468 ; 
      LAYER V1 ; 
        RECT 0.072 0.396 0.144 0.468 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.252 0.576 0.44 ; 
        RECT 0.424 0.252 0.576 0.324 ; 
      LAYER M2 ; 
        RECT 0.388 0.252 0.644 0.324 ; 
      LAYER V1 ; 
        RECT 0.452 0.252 0.524 0.324 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.252 0.868 0.324 ; 
        RECT 0.64 0.54 0.792 0.612 ; 
        RECT 0.72 0.252 0.792 0.612 ; 
      LAYER M2 ; 
        RECT 0.628 0.396 0.884 0.468 ; 
      LAYER V1 ; 
        RECT 0.72 0.396 0.792 0.468 ; 
    END 
  END C 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.252 0.108 0.9 0.18 ; 
        RECT 0.252 0.54 0.488 0.612 ; 
        RECT 0.252 0.108 0.324 0.612 ; 
      LAYER M2 ; 
        RECT 0.198 0.54 0.48 0.612 ; 
      LAYER V1 ; 
        RECT 0.312 0.54 0.384 0.612 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.828 0.684 1.352 0.756 ; 
      RECT 0.16 0.684 0.704 0.756 ; 
  END 
END AOI221xp25_ASAP7_6t_SL 


MACRO AOI221xp5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI221xp5_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.016 0.252 1.168 0.324 ; 
        RECT 1.016 0.54 1.164 0.612 ; 
        RECT 1.016 0.252 1.088 0.612 ; 
        RECT 0.924 0.384 1.088 0.456 ; 
      LAYER M2 ; 
        RECT 0.712 0.252 1.128 0.324 ; 
      LAYER V1 ; 
        RECT 1.036 0.252 1.108 0.324 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.292 0.464 1.448 0.612 ; 
        RECT 1.376 0.108 1.448 0.612 ; 
        RECT 1.236 0.108 1.448 0.18 ; 
      LAYER M2 ; 
        RECT 1.032 0.396 1.448 0.468 ; 
      LAYER V1 ; 
        RECT 1.376 0.396 1.448 0.468 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.212 0.188 0.36 ; 
        RECT 0.072 0.212 0.144 0.488 ; 
      LAYER M2 ; 
        RECT 0.096 0.252 0.512 0.324 ; 
      LAYER V1 ; 
        RECT 0.116 0.252 0.188 0.324 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.516 0.252 0.588 0.476 ; 
        RECT 0.432 0.252 0.588 0.324 ; 
      LAYER M2 ; 
        RECT 0.18 0.396 0.588 0.468 ; 
      LAYER V1 ; 
        RECT 0.516 0.396 0.588 0.468 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.636 0.54 0.892 0.612 ; 
        RECT 0.688 0.252 0.856 0.324 ; 
        RECT 0.72 0.252 0.792 0.612 ; 
      LAYER M2 ; 
        RECT 0.676 0.54 1.092 0.612 ; 
      LAYER V1 ; 
        RECT 0.696 0.54 0.768 0.612 ; 
    END 
  END C 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.26 0.108 0.9 0.18 ; 
        RECT 0.26 0.54 0.448 0.612 ; 
        RECT 0.26 0.108 0.332 0.612 ; 
      LAYER M2 ; 
        RECT 0.188 0.108 0.816 0.18 ; 
      LAYER V1 ; 
        RECT 0.396 0.108 0.468 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.808 0.684 1.352 0.756 ; 
      RECT 0.16 0.684 0.684 0.756 ; 
  END 
END AOI221xp5_ASAP7_6t_SL 


MACRO AOI222xp25_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI222xp25_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.232 0.144 0.584 ; 
      LAYER M2 ; 
        RECT 0.072 0.396 0.352 0.468 ; 
      LAYER V1 ; 
        RECT 0.072 0.396 0.144 0.468 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.252 0.576 0.468 ; 
        RECT 0.424 0.252 0.576 0.324 ; 
      LAYER M2 ; 
        RECT 0.412 0.252 0.748 0.324 ; 
      LAYER V1 ; 
        RECT 0.448 0.252 0.52 0.324 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.14 0.396 1.42 0.468 ; 
        RECT 1.348 0.252 1.42 0.468 ; 
        RECT 1.2 0.252 1.42 0.324 ; 
      LAYER M2 ; 
        RECT 1.148 0.252 1.484 0.324 ; 
      LAYER V1 ; 
        RECT 1.252 0.252 1.324 0.324 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.728 0.396 0.948 0.468 ; 
        RECT 0.728 0.252 0.948 0.324 ; 
        RECT 0.728 0.252 0.8 0.468 ; 
      LAYER M2 ; 
        RECT 0.656 0.396 0.952 0.468 ; 
      LAYER V1 ; 
        RECT 0.8 0.396 0.872 0.468 ; 
    END 
  END B2 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.664 0.464 1.812 0.612 ; 
        RECT 1.664 0.108 1.812 0.256 ; 
        RECT 1.664 0.108 1.736 0.612 ; 
        RECT 1.572 0.388 1.736 0.46 ; 
      LAYER M2 ; 
        RECT 1.444 0.396 1.84 0.468 ; 
      LAYER V1 ; 
        RECT 1.664 0.396 1.736 0.468 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.884 0.6 2.096 0.756 ; 
        RECT 2.024 0.108 2.096 0.756 ; 
        RECT 1.888 0.108 2.096 0.256 ; 
      LAYER M2 ; 
        RECT 1.788 0.684 2.096 0.756 ; 
      LAYER V1 ; 
        RECT 1.908 0.684 1.98 0.756 ; 
    END 
  END C2 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.252 0.108 1.352 0.18 ; 
        RECT 0.252 0.54 0.468 0.612 ; 
        RECT 0.252 0.108 0.324 0.612 ; 
      LAYER M2 ; 
        RECT 0.22 0.54 0.528 0.612 ; 
      LAYER V1 ; 
        RECT 0.328 0.54 0.4 0.612 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.368 0.684 1.784 0.756 ; 
      RECT 1.368 0.54 1.44 0.756 ; 
      RECT 0.796 0.54 1.44 0.612 ; 
      RECT 0.16 0.684 1.136 0.756 ; 
  END 
END AOI222xp25_ASAP7_6t_SL 


MACRO AOI22xp25_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI22xp25_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.124 0.464 0.272 0.612 ; 
        RECT 0.124 0.108 0.272 0.256 ; 
        RECT 0.124 0.108 0.196 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.42 0.392 0.564 0.464 ; 
        RECT 0.344 0.464 0.492 0.612 ; 
        RECT 0.42 0.108 0.492 0.612 ; 
        RECT 0.344 0.108 0.492 0.256 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.464 1.176 0.612 ; 
        RECT 1.104 0.108 1.176 0.612 ; 
        RECT 1.024 0.108 1.176 0.18 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.54 0.764 0.612 ; 
        RECT 0.692 0.108 0.764 0.612 ; 
        RECT 0.564 0.108 0.764 0.256 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.844 0.22 0.916 0.632 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.992 0.684 1.14 0.756 ; 
      RECT 0.16 0.684 0.704 0.756 ; 
    LAYER M2 ; 
      RECT 0.592 0.684 1.136 0.756 ; 
    LAYER V1 ; 
      RECT 1.044 0.684 1.116 0.756 ; 
      RECT 0.612 0.684 0.684 0.756 ; 
  END 
END AOI22xp25_ASAP7_6t_SL 


MACRO AOI22xp5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI22xp5_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.124 0.464 0.272 0.612 ; 
        RECT 0.124 0.108 0.272 0.256 ; 
        RECT 0.124 0.108 0.196 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.42 0.392 0.564 0.464 ; 
        RECT 0.344 0.464 0.492 0.612 ; 
        RECT 0.42 0.108 0.492 0.612 ; 
        RECT 0.344 0.108 0.492 0.256 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.464 1.176 0.612 ; 
        RECT 1.104 0.108 1.176 0.612 ; 
        RECT 1.024 0.108 1.176 0.18 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.54 0.764 0.612 ; 
        RECT 0.692 0.108 0.764 0.612 ; 
        RECT 0.564 0.108 0.764 0.256 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.844 0.22 0.916 0.632 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.992 0.684 1.14 0.756 ; 
      RECT 0.16 0.684 0.704 0.756 ; 
    LAYER M2 ; 
      RECT 0.592 0.684 1.136 0.756 ; 
    LAYER V1 ; 
      RECT 1.044 0.684 1.116 0.756 ; 
      RECT 0.612 0.684 0.684 0.756 ; 
  END 
END AOI22xp5_ASAP7_6t_SL 


MACRO AOI311xp33_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI311xp33_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.68 0.252 0.828 0.324 ; 
        RECT 0.72 0.252 0.792 0.488 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.54 0.576 0.612 ; 
        RECT 0.504 0.108 0.576 0.612 ; 
        RECT 0.376 0.108 0.576 0.18 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.36 0.468 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A3 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.86 0.54 1.008 0.612 ; 
        RECT 0.936 0.376 1.008 0.612 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.108 0.54 1.268 0.612 ; 
        RECT 1.12 0.252 1.268 0.324 ; 
        RECT 1.152 0.252 1.224 0.612 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.208 0.684 1.44 0.756 ; 
        RECT 1.368 0.108 1.44 0.756 ; 
        RECT 0.792 0.108 1.44 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.684 0.936 0.756 ; 
  END 
END AOI311xp33_ASAP7_6t_SL 


MACRO AOI31xp33_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI31xp33_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.636 0.464 0.816 0.612 ; 
        RECT 0.708 0.256 0.78 0.612 ; 
        RECT 0.664 0.256 0.78 0.328 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.464 0.564 0.612 ; 
        RECT 0.492 0.108 0.564 0.612 ; 
        RECT 0.364 0.108 0.564 0.256 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.068 0.608 0.276 0.756 ; 
        RECT 0.068 0.108 0.272 0.256 ; 
        RECT 0.068 0.108 0.14 0.756 ; 
    END 
  END A3 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.908 0.252 1.06 0.332 ; 
        RECT 0.9 0.464 1.048 0.612 ; 
        RECT 0.936 0.252 1.008 0.612 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.16 0.108 1.232 0.728 ; 
        RECT 0.808 0.108 1.232 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.684 0.92 0.756 ; 
  END 
END AOI31xp33_ASAP7_6t_SL 


MACRO AOI31xp67_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI31xp67_ASAP7_6t_SL 0 0 ; 
  SIZE 2.808 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.052 0.396 2.756 0.468 ; 
        RECT 2.684 0.252 2.756 0.468 ; 
        RECT 2.536 0.252 2.756 0.324 ; 
        RECT 2.32 0.684 2.468 0.756 ; 
        RECT 2.32 0.396 2.392 0.756 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.092 0.396 1.864 0.468 ; 
        RECT 1.092 0.54 1.312 0.612 ; 
        RECT 1.092 0.108 1.312 0.18 ; 
        RECT 1.092 0.108 1.164 0.612 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.38 0.468 ; 
        RECT 0.072 0.54 0.292 0.612 ; 
        RECT 0.072 0.108 0.252 0.18 ; 
        RECT 0.072 0.108 0.144 0.612 ; 
    END 
  END A3 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.616 0.392 0.836 0.464 ; 
        RECT 0.484 0.54 0.688 0.612 ; 
        RECT 0.616 0.252 0.688 0.612 ; 
        RECT 0.468 0.252 0.688 0.324 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.808 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.808 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.828 0.54 2.652 0.612 ; 
      LAYER M1 ; 
        RECT 2.516 0.54 2.696 0.612 ; 
        RECT 0.8 0.54 1.02 0.612 ; 
        RECT 0.948 0.108 1.02 0.612 ; 
        RECT 0.808 0.108 1.02 0.18 ; 
      LAYER V1 ; 
        RECT 0.928 0.54 1 0.612 ; 
        RECT 2.56 0.54 2.632 0.612 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 2.104 0.108 2.652 0.18 ; 
      RECT 1.456 0.252 2.412 0.324 ; 
      RECT 0.16 0.684 2.216 0.756 ; 
      RECT 1.632 0.108 1.788 0.18 ; 
      RECT 0.376 0.108 0.524 0.18 ; 
    LAYER M2 ; 
      RECT 0.376 0.108 1.788 0.18 ; 
    LAYER V1 ; 
      RECT 1.692 0.108 1.764 0.18 ; 
      RECT 0.396 0.108 0.468 0.18 ; 
  END 
END AOI31xp67_ASAP7_6t_SL 


MACRO AOI321xp17_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI321xp17_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.488 ; 
      LAYER M2 ; 
        RECT 0.632 0.396 0.888 0.468 ; 
      LAYER V1 ; 
        RECT 0.72 0.396 0.792 0.468 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.54 0.576 0.612 ; 
        RECT 0.504 0.108 0.576 0.612 ; 
        RECT 0.376 0.108 0.576 0.18 ; 
      LAYER M2 ; 
        RECT 0.388 0.54 0.652 0.612 ; 
      LAYER V1 ; 
        RECT 0.496 0.54 0.568 0.612 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
      LAYER M2 ; 
        RECT 0.072 0.396 0.424 0.468 ; 
      LAYER V1 ; 
        RECT 0.072 0.396 0.144 0.468 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.108 0.108 1.268 0.18 ; 
        RECT 1.14 0.108 1.212 0.476 ; 
      LAYER M2 ; 
        RECT 1.028 0.396 1.284 0.468 ; 
      LAYER V1 ; 
        RECT 1.14 0.396 1.212 0.468 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.44 0.252 1.512 0.44 ; 
        RECT 1.364 0.252 1.512 0.324 ; 
      LAYER M2 ; 
        RECT 1.356 0.252 1.612 0.324 ; 
      LAYER V1 ; 
        RECT 1.404 0.252 1.476 0.324 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.54 1.084 0.612 ; 
        RECT 0.936 0.28 1.008 0.612 ; 
      LAYER M2 ; 
        RECT 0.848 0.54 1.112 0.612 ; 
      LAYER V1 ; 
        RECT 0.944 0.54 1.016 0.612 ; 
    END 
  END C 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.26 0.54 1.656 0.612 ; 
        RECT 1.584 0.108 1.656 0.612 ; 
        RECT 1.424 0.108 1.656 0.18 ; 
        RECT 0.792 0.108 0.952 0.18 ; 
      LAYER M2 ; 
        RECT 0.828 0.108 1.568 0.18 ; 
      LAYER V1 ; 
        RECT 0.828 0.108 0.9 0.18 ; 
        RECT 1.476 0.108 1.548 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.024 0.684 1.584 0.756 ; 
      RECT 0.376 0.684 0.9 0.756 ; 
  END 
END AOI321xp17_ASAP7_6t_SL 


MACRO AOI322xp17_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI322xp17_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.54 0.284 0.612 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.612 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.564 0.396 0.88 0.468 ; 
      LAYER M1 ; 
        RECT 0.636 0.396 0.784 0.468 ; 
        RECT 0.636 0.244 0.708 0.468 ; 
      LAYER V1 ; 
        RECT 0.68 0.396 0.752 0.468 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.808 0.252 1.08 0.324 ; 
      LAYER M1 ; 
        RECT 0.936 0.252 1.008 0.44 ; 
        RECT 0.82 0.252 1.008 0.324 ; 
      LAYER V1 ; 
        RECT 0.828 0.252 0.9 0.324 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 1.084 0.54 1.448 0.612 ; 
      LAYER M1 ; 
        RECT 1.168 0.54 1.332 0.612 ; 
        RECT 1.12 0.108 1.268 0.18 ; 
        RECT 1.168 0.352 1.24 0.612 ; 
        RECT 1.152 0.108 1.224 0.424 ; 
      LAYER V1 ; 
        RECT 1.208 0.54 1.28 0.612 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.304 0.252 0.612 0.324 ; 
      LAYER M1 ; 
        RECT 0.336 0.396 0.564 0.468 ; 
        RECT 0.492 0.108 0.564 0.468 ; 
        RECT 0.376 0.108 0.564 0.18 ; 
      LAYER V1 ; 
        RECT 0.492 0.252 0.564 0.324 ; 
    END 
  END B1 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 1.512 0.252 1.792 0.324 ; 
      LAYER M1 ; 
        RECT 1.648 0.252 1.72 0.44 ; 
        RECT 1.552 0.252 1.72 0.324 ; 
      LAYER V1 ; 
        RECT 1.56 0.252 1.632 0.324 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 1.304 0.396 1.6 0.468 ; 
      LAYER M1 ; 
        RECT 1.368 0.396 1.516 0.468 ; 
        RECT 1.368 0.108 1.516 0.18 ; 
        RECT 1.368 0.108 1.44 0.468 ; 
      LAYER V1 ; 
        RECT 1.404 0.396 1.476 0.468 ; 
    END 
  END C2 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.808 0.108 1.784 0.18 ; 
      LAYER M1 ; 
        RECT 1.456 0.54 1.872 0.612 ; 
        RECT 1.8 0.108 1.872 0.612 ; 
        RECT 1.652 0.108 1.872 0.18 ; 
        RECT 0.776 0.108 0.996 0.18 ; 
      LAYER V1 ; 
        RECT 0.828 0.108 0.9 0.18 ; 
        RECT 1.692 0.108 1.764 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.684 0.704 0.756 ; 
      RECT 0.408 0.54 0.48 0.756 ; 
      RECT 0.408 0.54 1.068 0.612 ; 
      RECT 0.828 0.684 1.8 0.756 ; 
  END 
END AOI322xp17_ASAP7_6t_SL 


MACRO AOI32xp33_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI32xp33_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.064 0.108 0.272 0.18 ; 
        RECT 0.064 0.108 0.136 0.508 ; 
      LAYER M2 ; 
        RECT 0.152 0.108 0.672 0.18 ; 
      LAYER V1 ; 
        RECT 0.18 0.108 0.252 0.18 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.312 0.396 0.596 0.468 ; 
      LAYER M2 ; 
        RECT 0.244 0.396 0.652 0.468 ; 
      LAYER V1 ; 
        RECT 0.4 0.396 0.472 0.468 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.672 0.54 0.884 0.612 ; 
        RECT 0.72 0.352 0.792 0.612 ; 
      LAYER M2 ; 
        RECT 0.588 0.54 0.996 0.612 ; 
      LAYER V1 ; 
        RECT 0.772 0.54 0.844 0.612 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.928 0.252 1.08 0.324 ; 
        RECT 0.928 0.252 1 0.472 ; 
      LAYER M2 ; 
        RECT 0.86 0.252 1.228 0.324 ; 
      LAYER V1 ; 
        RECT 0.996 0.252 1.068 0.324 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.116 0.396 1.308 0.468 ; 
        RECT 1.236 0.28 1.308 0.468 ; 
      LAYER M2 ; 
        RECT 0.972 0.396 1.38 0.468 ; 
      LAYER V1 ; 
        RECT 1.136 0.396 1.208 0.468 ; 
    END 
  END B2 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.044 0.54 1.452 0.612 ; 
        RECT 1.38 0.108 1.452 0.612 ; 
        RECT 0.592 0.108 1.452 0.18 ; 
        RECT 1.044 0.54 1.116 0.704 ; 
      LAYER M2 ; 
        RECT 0.836 0.108 1.352 0.18 ; 
      LAYER V1 ; 
        RECT 1.26 0.108 1.332 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.24 0.684 1.388 0.756 ; 
      RECT 0.376 0.684 0.92 0.756 ; 
    LAYER M2 ; 
      RECT 0.592 0.684 1.352 0.756 ; 
    LAYER V1 ; 
      RECT 1.26 0.684 1.332 0.756 ; 
      RECT 0.612 0.684 0.684 0.756 ; 
  END 
END AOI32xp33_ASAP7_6t_SL 


MACRO AOI331xp17_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI331xp17_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.54 0.896 0.612 ; 
        RECT 0.72 0.28 0.792 0.612 ; 
      LAYER M2 ; 
        RECT 0.728 0.54 1.088 0.612 ; 
      LAYER V1 ; 
        RECT 0.8 0.54 0.872 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.54 0.62 0.612 ; 
        RECT 0.376 0.108 0.62 0.18 ; 
        RECT 0.504 0.108 0.576 0.612 ; 
      LAYER M2 ; 
        RECT 0.354 0.252 0.71 0.324 ; 
      LAYER V1 ; 
        RECT 0.504 0.252 0.576 0.324 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.684 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
      LAYER M2 ; 
        RECT 0.152 0.684 0.544 0.756 ; 
      LAYER V1 ; 
        RECT 0.18 0.684 0.252 0.756 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.396 1.084 0.468 ; 
        RECT 0.936 0.28 1.008 0.468 ; 
      LAYER M2 ; 
        RECT 0.688 0.396 1.192 0.468 ; 
      LAYER V1 ; 
        RECT 0.948 0.396 1.02 0.468 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.112 0.108 1.26 0.18 ; 
        RECT 1.152 0.108 1.224 0.352 ; 
      LAYER M2 ; 
        RECT 0.848 0.252 1.244 0.324 ; 
      LAYER V1 ; 
        RECT 1.152 0.252 1.224 0.324 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.108 1.516 0.18 ; 
        RECT 1.368 0.108 1.44 0.432 ; 
      LAYER M2 ; 
        RECT 1.368 0.252 1.68 0.324 ; 
      LAYER V1 ; 
        RECT 1.368 0.252 1.44 0.324 ; 
    END 
  END B3 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.648 0.28 1.72 0.56 ; 
      LAYER M2 ; 
        RECT 1.456 0.396 1.812 0.468 ; 
      LAYER V1 ; 
        RECT 1.648 0.396 1.72 0.468 ; 
    END 
  END C 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.672 0.684 1.872 0.756 ; 
        RECT 1.8 0.108 1.872 0.756 ; 
        RECT 1.64 0.108 1.872 0.18 ; 
        RECT 0.78 0.108 0.948 0.18 ; 
      LAYER M2 ; 
        RECT 0.804 0.108 1.804 0.18 ; 
      LAYER V1 ; 
        RECT 0.828 0.108 0.9 0.18 ; 
        RECT 1.692 0.108 1.764 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.476 0.54 1.548 0.724 ; 
      RECT 1.024 0.54 1.548 0.612 ; 
      RECT 0.396 0.684 1.352 0.756 ; 
  END 
END AOI331xp17_ASAP7_6t_SL 


MACRO AOI332xp17_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI332xp17_ASAP7_6t_SL 0 0 ; 
  SIZE 2.376 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.636 0.388 0.804 0.46 ; 
        RECT 0.636 0.108 0.708 0.632 ; 
        RECT 0.376 0.108 0.708 0.18 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.54 0.564 0.612 ; 
        RECT 0.492 0.252 0.564 0.612 ; 
        RECT 0.32 0.252 0.564 0.324 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.252 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.828 0.54 0.996 0.612 ; 
        RECT 0.924 0.108 0.996 0.612 ; 
        RECT 0.808 0.108 0.996 0.18 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.068 0.108 1.332 0.18 ; 
        RECT 1.068 0.396 1.288 0.468 ; 
        RECT 1.068 0.108 1.14 0.468 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.428 0.396 1.664 0.468 ; 
        RECT 1.24 0.252 1.648 0.324 ; 
        RECT 1.428 0.252 1.5 0.468 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.228 0.204 2.3 0.56 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.792 0.396 2.012 0.468 ; 
        RECT 1.94 0.252 2.012 0.468 ; 
        RECT 1.78 0.252 2.012 0.324 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.376 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.928 0.54 2.156 0.612 ; 
        RECT 2.084 0.108 2.156 0.612 ; 
        RECT 1.456 0.108 2.156 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.732 0.684 2.272 0.756 ; 
      RECT 1.732 0.54 1.804 0.756 ; 
      RECT 1.1 0.54 1.804 0.612 ; 
      RECT 0.804 0.684 1.568 0.756 ; 
      RECT 0.376 0.684 0.54 0.756 ; 
    LAYER M2 ; 
      RECT 0.396 0.684 0.936 0.756 ; 
    LAYER V1 ; 
      RECT 0.828 0.684 0.9 0.756 ; 
      RECT 0.396 0.684 0.468 0.756 ; 
  END 
END AOI332xp17_ASAP7_6t_SL 


MACRO AOI333xp17_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI333xp17_ASAP7_6t_SL 0 0 ; 
  SIZE 2.808 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.32 0.108 2.648 0.18 ; 
        RECT 2.552 0.108 2.624 0.516 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.236 0.396 2.468 0.468 ; 
        RECT 2.396 0.252 2.468 0.468 ; 
        RECT 2.236 0.252 2.468 0.324 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.856 0.396 2.088 0.468 ; 
        RECT 1.856 0.252 2.084 0.324 ; 
        RECT 1.856 0.252 1.928 0.468 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.108 1.136 0.18 ; 
        RECT 0.948 0.108 1.02 0.464 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.164 0.396 1.44 0.468 ; 
        RECT 1.368 0.252 1.44 0.468 ; 
        RECT 1.18 0.252 1.44 0.324 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.556 0.396 1.784 0.468 ; 
        RECT 1.712 0.252 1.784 0.468 ; 
        RECT 1.564 0.252 1.784 0.324 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.712 0.54 0.92 0.612 ; 
        RECT 0.712 0.268 0.784 0.612 ; 
        RECT 0.636 0.268 0.784 0.352 ; 
        RECT 0.636 0.108 0.708 0.352 ; 
        RECT 0.42 0.108 0.708 0.18 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.344 0.54 0.564 0.612 ; 
        RECT 0.492 0.252 0.564 0.612 ; 
        RECT 0.32 0.252 0.564 0.324 ; 
    END 
  END C2 
  PIN C3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 0.28 0.18 ; 
        RECT 0.072 0.108 0.144 0.652 ; 
    END 
  END C3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.808 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.808 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 2.084 0.684 2.72 0.756 ; 
      LAYER M1 ; 
        RECT 2.532 0.684 2.768 0.756 ; 
        RECT 2.696 0.256 2.768 0.756 ; 
        RECT 2.02 0.684 2.216 0.756 ; 
      LAYER V1 ; 
        RECT 2.124 0.684 2.196 0.756 ; 
        RECT 2.556 0.684 2.628 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 2.34 0.54 2.412 0.704 ; 
      RECT 1.06 0.54 1.132 0.704 ; 
      RECT 1.06 0.54 2.412 0.612 ; 
      RECT 1.26 0.108 2.196 0.18 ; 
      RECT 1.26 0.684 1.572 0.756 ; 
      RECT 0.748 0.684 0.92 0.756 ; 
      RECT 0.344 0.684 0.54 0.756 ; 
    LAYER M2 ; 
      RECT 0.376 0.684 1.572 0.756 ; 
    LAYER V1 ; 
      RECT 1.476 0.684 1.548 0.756 ; 
      RECT 0.828 0.684 0.9 0.756 ; 
      RECT 0.396 0.684 0.468 0.756 ; 
  END 
END AOI333xp17_ASAP7_6t_SL 


MACRO AOI33xp33_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI33xp33_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.684 0.22 0.756 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.344 0.396 0.568 0.468 ; 
        RECT 0.344 0.108 0.492 0.18 ; 
        RECT 0.26 0.54 0.416 0.612 ; 
        RECT 0.344 0.108 0.416 0.612 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.644 0.54 0.792 0.612 ; 
        RECT 0.72 0.252 0.792 0.612 ; 
        RECT 0.536 0.252 0.792 0.324 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.008 0.108 1.248 0.18 ; 
        RECT 1.008 0.396 1.156 0.468 ; 
        RECT 1.008 0.108 1.08 0.468 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.284 0.396 1.524 0.468 ; 
        RECT 1.452 0.108 1.524 0.468 ; 
        RECT 1.376 0.108 1.524 0.18 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.836 0.108 1.908 0.66 ; 
        RECT 1.648 0.396 1.908 0.468 ; 
        RECT 1.76 0.108 1.908 0.18 ; 
    END 
  END B3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.692 0.54 1.764 0.704 ; 
        RECT 0.864 0.54 1.764 0.612 ; 
        RECT 0.864 0.108 0.936 0.612 ; 
        RECT 0.704 0.108 0.936 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.344 0.684 1.568 0.756 ; 
  END 
END AOI33xp33_ASAP7_6t_SL 


MACRO BUFx10_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx10_ASAP7_6t_SL 0 0 ; 
  SIZE 3.024 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.38 0.468 ; 
        RECT 0.072 0.684 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.024 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.024 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.684 2.952 0.756 ; 
        RECT 2.88 0.108 2.952 0.756 ; 
        RECT 0.808 0.108 2.952 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.396 0.684 0.576 0.756 ; 
      RECT 0.504 0.108 0.576 0.756 ; 
      RECT 0.504 0.396 2.756 0.468 ; 
      RECT 0.396 0.108 0.576 0.18 ; 
  END 
END BUFx10_ASAP7_6t_SL 


MACRO BUFx12_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx12_ASAP7_6t_SL 0 0 ; 
  SIZE 3.456 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.456 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.456 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.684 3.384 0.756 ; 
        RECT 3.312 0.108 3.384 0.756 ; 
        RECT 0.808 0.108 3.384 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.684 0.576 0.756 ; 
      RECT 0.504 0.108 0.576 0.756 ; 
      RECT 0.504 0.396 3.188 0.468 ; 
      RECT 0.376 0.108 0.576 0.18 ; 
  END 
END BUFx12_ASAP7_6t_SL 


MACRO BUFx12q_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx12q_ASAP7_6t_SL 0 0 ; 
  SIZE 3.888 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.08 0.396 0.38 0.468 ; 
        RECT 0.08 0.608 0.272 0.756 ; 
        RECT 0.08 0.108 0.272 0.256 ; 
        RECT 0.08 0.108 0.152 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.888 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.888 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.24 0.684 3.816 0.756 ; 
        RECT 3.744 0.108 3.816 0.756 ; 
        RECT 1.24 0.108 3.816 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.684 1.116 0.756 ; 
      RECT 1.044 0.108 1.116 0.756 ; 
      RECT 1.044 0.396 1.244 0.468 ; 
      RECT 0.376 0.108 1.116 0.18 ; 
  END 
END BUFx12q_ASAP7_6t_SL 


MACRO BUFx16q_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx16q_ASAP7_6t_SL 0 0 ; 
  SIZE 4.752 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.068 0.396 0.38 0.468 ; 
        RECT 0.068 0.608 0.272 0.756 ; 
        RECT 0.068 0.108 0.272 0.256 ; 
        RECT 0.068 0.108 0.14 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 4.752 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.752 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.24 0.684 4.68 0.756 ; 
        RECT 4.608 0.108 4.68 0.756 ; 
        RECT 1.24 0.108 4.68 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.684 1.008 0.756 ; 
      RECT 0.936 0.108 1.008 0.756 ; 
      RECT 0.936 0.396 4.484 0.468 ; 
      RECT 0.376 0.108 1.008 0.18 ; 
  END 
END BUFx16q_ASAP7_6t_SL 


MACRO BUFx24_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx24_ASAP7_6t_SL 0 0 ; 
  SIZE 6.48 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.744 0.468 ; 
        RECT 0.072 0.684 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 6.48 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 6.48 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.24 0.684 6.408 0.756 ; 
        RECT 6.336 0.108 6.408 0.756 ; 
        RECT 1.24 0.108 6.408 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.396 0.684 1.008 0.756 ; 
      RECT 0.936 0.108 1.008 0.756 ; 
      RECT 0.936 0.396 6.212 0.468 ; 
      RECT 0.396 0.108 1.008 0.18 ; 
  END 
END BUFx24_ASAP7_6t_SL 


MACRO BUFx2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx2_ASAP7_6t_SL 0 0 ; 
  SIZE 1.08 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.312 0.468 ; 
        RECT 0.072 0.54 0.292 0.612 ; 
        RECT 0.072 0.252 0.292 0.324 ; 
        RECT 0.072 0.252 0.144 0.612 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.08 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.08 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.684 1.008 0.756 ; 
        RECT 0.936 0.108 1.008 0.756 ; 
        RECT 0.592 0.108 1.008 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.684 0.488 0.756 ; 
      RECT 0.416 0.108 0.488 0.756 ; 
      RECT 0.416 0.396 0.812 0.468 ; 
      RECT 0.16 0.108 0.488 0.18 ; 
  END 
END BUFx2_ASAP7_6t_SL 


MACRO BUFx3_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx3_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.04 0.396 0.312 0.468 ; 
        RECT 0.04 0.54 0.296 0.612 ; 
        RECT 0.04 0.252 0.296 0.324 ; 
        RECT 0.04 0.252 0.112 0.612 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.684 1.224 0.756 ; 
        RECT 1.152 0.108 1.224 0.756 ; 
        RECT 0.592 0.108 1.224 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.684 0.488 0.756 ; 
      RECT 0.416 0.108 0.488 0.756 ; 
      RECT 0.416 0.396 1.028 0.468 ; 
      RECT 0.16 0.108 0.488 0.18 ; 
  END 
END BUFx3_ASAP7_6t_SL 


MACRO BUFx4_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx4_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.04 0.396 0.312 0.468 ; 
        RECT 0.04 0.54 0.272 0.612 ; 
        RECT 0.04 0.252 0.272 0.324 ; 
        RECT 0.04 0.252 0.112 0.612 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.684 1.428 0.756 ; 
        RECT 1.356 0.108 1.428 0.756 ; 
        RECT 0.592 0.108 1.428 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.684 0.488 0.756 ; 
      RECT 0.416 0.108 0.488 0.756 ; 
      RECT 0.416 0.396 1.244 0.468 ; 
      RECT 0.16 0.108 0.488 0.18 ; 
  END 
END BUFx4_ASAP7_6t_SL 


MACRO BUFx4q_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx4q_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.496 0.468 ; 
        RECT 0.072 0.684 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.684 1.648 0.756 ; 
        RECT 1.576 0.108 1.648 0.756 ; 
        RECT 0.808 0.108 1.648 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.396 0.684 0.708 0.756 ; 
      RECT 0.636 0.108 0.708 0.756 ; 
      RECT 0.636 0.396 1.46 0.468 ; 
      RECT 0.396 0.108 0.708 0.18 ; 
  END 
END BUFx4q_ASAP7_6t_SL 


MACRO BUFx5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx5_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.044 0.396 0.312 0.468 ; 
        RECT 0.044 0.54 0.264 0.612 ; 
        RECT 0.044 0.252 0.264 0.324 ; 
        RECT 0.044 0.252 0.116 0.612 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.684 1.656 0.756 ; 
        RECT 1.584 0.108 1.656 0.756 ; 
        RECT 0.592 0.108 1.656 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.684 0.488 0.756 ; 
      RECT 0.416 0.108 0.488 0.756 ; 
      RECT 0.416 0.396 1.46 0.468 ; 
      RECT 0.16 0.108 0.488 0.18 ; 
  END 
END BUFx5_ASAP7_6t_SL 


MACRO BUFx6q_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx6q_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.336 0.468 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.684 2.088 0.756 ; 
        RECT 2.016 0.108 2.088 0.756 ; 
        RECT 0.808 0.108 2.088 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.684 0.576 0.756 ; 
      RECT 0.504 0.108 0.576 0.756 ; 
      RECT 0.504 0.396 1.892 0.468 ; 
      RECT 0.376 0.108 0.576 0.18 ; 
  END 
END BUFx6q_ASAP7_6t_SL 


MACRO BUFx8_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx8_ASAP7_6t_SL 0 0 ; 
  SIZE 2.592 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.38 0.468 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.592 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.684 2.52 0.756 ; 
        RECT 2.448 0.108 2.52 0.756 ; 
        RECT 0.808 0.108 2.52 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.684 0.576 0.756 ; 
      RECT 0.504 0.108 0.576 0.756 ; 
      RECT 0.504 0.396 2.324 0.468 ; 
      RECT 0.376 0.108 0.576 0.18 ; 
  END 
END BUFx8_ASAP7_6t_SL 


MACRO CKINVDCx10_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN CKINVDCx10_ASAP7_6t_SL 0 0 ; 
  SIZE 5.184 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.284 0.396 4.68 0.468 ; 
        RECT 4.48 0.108 4.552 0.468 ; 
        RECT 0.072 0.108 4.552 0.18 ; 
        RECT 2.988 0.396 3.256 0.468 ; 
        RECT 3.184 0.108 3.256 0.468 ; 
        RECT 1.496 0.396 1.764 0.468 ; 
        RECT 1.496 0.108 1.568 0.468 ; 
        RECT 0.072 0.396 0.468 0.468 ; 
        RECT 0.072 0.684 0.272 0.756 ; 
        RECT 0.072 0.108 0.148 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 5.184 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.184 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.684 4.896 0.756 ; 
        RECT 4.824 0.108 4.896 0.756 ; 
        RECT 4.696 0.108 4.896 0.18 ; 
        RECT 4.112 0.252 4.376 0.324 ; 
        RECT 4.112 0.252 4.184 0.756 ; 
        RECT 2.816 0.252 3.08 0.324 ; 
        RECT 2.816 0.252 2.888 0.756 ; 
        RECT 1.864 0.252 1.936 0.756 ; 
        RECT 1.672 0.252 1.936 0.324 ; 
        RECT 0.568 0.252 0.64 0.756 ; 
        RECT 0.376 0.252 0.64 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 3.744 0.396 3.968 0.468 ; 
      RECT 3.744 0.252 3.816 0.468 ; 
      RECT 3.4 0.252 4.008 0.324 ; 
      RECT 3.324 0.54 3.944 0.612 ; 
      RECT 3.528 0.396 3.6 0.612 ; 
      RECT 3.368 0.396 3.6 0.468 ; 
      RECT 2.104 0.54 2.7 0.612 ; 
      RECT 2.448 0.396 2.52 0.612 ; 
      RECT 2.448 0.396 2.68 0.468 ; 
      RECT 2.08 0.396 2.304 0.468 ; 
      RECT 2.232 0.252 2.304 0.468 ; 
      RECT 2.04 0.252 2.648 0.324 ; 
      RECT 0.808 0.54 1.428 0.612 ; 
      RECT 1.152 0.396 1.224 0.612 ; 
      RECT 1.152 0.396 1.384 0.468 ; 
      RECT 0.784 0.396 1.008 0.468 ; 
      RECT 0.936 0.252 1.008 0.468 ; 
      RECT 0.744 0.252 1.352 0.324 ; 
  END 
END CKINVDCx10_ASAP7_6t_SL 


MACRO CKINVDCx11_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN CKINVDCx11_ASAP7_6t_SL 0 0 ; 
  SIZE 5.616 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.148 0.396 5.456 0.468 ; 
        RECT 5.344 0.108 5.456 0.468 ; 
        RECT 0.16 0.108 5.456 0.18 ; 
        RECT 3.42 0.396 3.924 0.468 ; 
        RECT 3.636 0.108 3.708 0.468 ; 
        RECT 1.692 0.396 2.196 0.468 ; 
        RECT 1.904 0.108 1.976 0.468 ; 
        RECT 0.16 0.396 0.468 0.468 ; 
        RECT 0.16 0.108 0.268 0.468 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 5.616 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.616 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.368 0.684 5.24 0.756 ; 
        RECT 4.976 0.252 5.22 0.324 ; 
        RECT 4.976 0.252 5.048 0.756 ; 
        RECT 4.024 0.252 4.096 0.756 ; 
        RECT 3.824 0.252 4.096 0.324 ; 
        RECT 3.232 0.252 3.492 0.324 ; 
        RECT 3.232 0.252 3.32 0.756 ; 
        RECT 2.3 0.252 2.372 0.756 ; 
        RECT 2.096 0.252 2.372 0.324 ; 
        RECT 1.52 0.252 1.764 0.324 ; 
        RECT 1.52 0.252 1.592 0.756 ; 
        RECT 0.568 0.252 0.64 0.756 ; 
        RECT 0.368 0.252 0.64 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 4.608 0.396 4.832 0.468 ; 
      RECT 4.608 0.252 4.68 0.468 ; 
      RECT 4.264 0.252 4.872 0.324 ; 
      RECT 4.216 0.54 4.808 0.612 ; 
      RECT 4.392 0.396 4.464 0.612 ; 
      RECT 4.232 0.396 4.464 0.468 ; 
      RECT 2.536 0.54 3.128 0.612 ; 
      RECT 2.88 0.396 2.952 0.612 ; 
      RECT 2.88 0.396 3.112 0.468 ; 
      RECT 2.512 0.396 2.736 0.468 ; 
      RECT 2.664 0.252 2.736 0.468 ; 
      RECT 2.472 0.252 3.08 0.324 ; 
      RECT 0.808 0.54 1.396 0.612 ; 
      RECT 1.152 0.396 1.224 0.612 ; 
      RECT 1.152 0.396 1.384 0.468 ; 
      RECT 0.784 0.396 1.008 0.468 ; 
      RECT 0.936 0.252 1.008 0.468 ; 
      RECT 0.744 0.252 1.352 0.324 ; 
  END 
END CKINVDCx11_ASAP7_6t_SL 


MACRO CKINVDCx12_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN CKINVDCx12_ASAP7_6t_SL 0 0 ; 
  SIZE 5.616 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.124 0.396 5.416 0.468 ; 
        RECT 5.344 0.108 5.416 0.468 ; 
        RECT 0.196 0.108 5.416 0.18 ; 
        RECT 3.4 0.396 3.944 0.468 ; 
        RECT 3.636 0.108 3.708 0.468 ; 
        RECT 1.672 0.396 2.216 0.468 ; 
        RECT 1.904 0.108 1.976 0.468 ; 
        RECT 0.196 0.396 0.488 0.468 ; 
        RECT 0.196 0.108 0.268 0.468 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 5.616 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.616 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.368 0.684 5.244 0.756 ; 
        RECT 4.948 0.252 5.24 0.324 ; 
        RECT 4.948 0.252 5.02 0.756 ; 
        RECT 4.044 0.252 4.116 0.756 ; 
        RECT 3.824 0.252 4.116 0.324 ; 
        RECT 3.212 0.252 3.512 0.324 ; 
        RECT 3.212 0.252 3.292 0.756 ; 
        RECT 2.332 0.252 2.412 0.756 ; 
        RECT 2.096 0.252 2.412 0.324 ; 
        RECT 1.488 0.252 1.784 0.324 ; 
        RECT 1.488 0.252 1.56 0.756 ; 
        RECT 0.608 0.252 0.68 0.756 ; 
        RECT 0.368 0.252 0.68 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 4.608 0.396 4.836 0.468 ; 
      RECT 4.608 0.252 4.68 0.468 ; 
      RECT 4.236 0.252 4.84 0.324 ; 
      RECT 4.236 0.54 4.808 0.612 ; 
      RECT 4.392 0.396 4.464 0.612 ; 
      RECT 4.236 0.396 4.464 0.468 ; 
      RECT 2.536 0.54 3.1 0.612 ; 
      RECT 2.88 0.396 2.952 0.612 ; 
      RECT 2.88 0.396 3.1 0.468 ; 
      RECT 2.512 0.396 2.736 0.468 ; 
      RECT 2.664 0.252 2.736 0.468 ; 
      RECT 2.512 0.252 3.08 0.324 ; 
      RECT 0.808 0.54 1.384 0.612 ; 
      RECT 1.152 0.396 1.224 0.612 ; 
      RECT 1.152 0.396 1.384 0.468 ; 
      RECT 0.784 0.396 1.008 0.468 ; 
      RECT 0.936 0.252 1.008 0.468 ; 
      RECT 0.784 0.252 1.352 0.324 ; 
  END 
END CKINVDCx12_ASAP7_6t_SL 


MACRO CKINVDCx14_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN CKINVDCx14_ASAP7_6t_SL 0 0 ; 
  SIZE 6.048 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.216 0.396 5.588 0.468 ; 
        RECT 5.364 0.108 5.436 0.468 ; 
        RECT 0.16 0.108 5.436 0.18 ; 
        RECT 3.488 0.396 3.856 0.468 ; 
        RECT 3.636 0.108 3.708 0.468 ; 
        RECT 1.756 0.396 2.124 0.468 ; 
        RECT 1.904 0.108 1.976 0.468 ; 
        RECT 0.16 0.396 0.404 0.468 ; 
        RECT 0.16 0.108 0.256 0.468 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 6.048 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 6.048 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 5.888 0.756 ; 
        RECT 5.816 0.108 5.888 0.756 ; 
        RECT 5.536 0.108 5.888 0.18 ; 
        RECT 5.04 0.252 5.26 0.324 ; 
        RECT 5.04 0.252 5.112 0.756 ; 
        RECT 3.96 0.252 4.032 0.756 ; 
        RECT 3.808 0.252 4.032 0.324 ; 
        RECT 3.312 0.252 3.532 0.324 ; 
        RECT 3.312 0.252 3.384 0.756 ; 
        RECT 2.232 0.252 2.304 0.756 ; 
        RECT 2.084 0.252 2.304 0.324 ; 
        RECT 1.584 0.252 1.804 0.324 ; 
        RECT 1.584 0.252 1.656 0.756 ; 
        RECT 0.504 0.252 0.576 0.756 ; 
        RECT 0.356 0.252 0.576 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 4.608 0.396 4.832 0.468 ; 
      RECT 4.608 0.252 4.68 0.468 ; 
      RECT 4.264 0.252 4.872 0.324 ; 
      RECT 4.188 0.54 4.808 0.612 ; 
      RECT 4.392 0.396 4.464 0.612 ; 
      RECT 4.232 0.396 4.464 0.468 ; 
      RECT 2.536 0.54 3.156 0.612 ; 
      RECT 2.88 0.396 2.952 0.612 ; 
      RECT 2.88 0.396 3.112 0.468 ; 
      RECT 2.512 0.396 2.736 0.468 ; 
      RECT 2.664 0.252 2.736 0.468 ; 
      RECT 2.472 0.252 3.08 0.324 ; 
      RECT 0.808 0.54 1.428 0.612 ; 
      RECT 1.152 0.396 1.224 0.612 ; 
      RECT 1.152 0.396 1.384 0.468 ; 
      RECT 0.784 0.396 1.008 0.468 ; 
      RECT 0.936 0.252 1.008 0.468 ; 
      RECT 0.744 0.252 1.352 0.324 ; 
  END 
END CKINVDCx14_ASAP7_6t_SL 


MACRO CKINVDCx16_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN CKINVDCx16_ASAP7_6t_SL 0 0 ; 
  SIZE 6.48 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 6.208 0.684 6.408 0.756 ; 
        RECT 6.336 0.108 6.408 0.756 ; 
        RECT 5.692 0.396 6.408 0.468 ; 
        RECT 0.608 0.108 6.408 0.18 ; 
        RECT 3.92 0.396 4.288 0.468 ; 
        RECT 4.068 0.108 4.14 0.468 ; 
        RECT 2.188 0.396 2.556 0.468 ; 
        RECT 2.336 0.108 2.408 0.468 ; 
        RECT 0.472 0.396 0.828 0.468 ; 
        RECT 0.608 0.108 0.68 0.468 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 6.48 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 6.48 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.228 0.684 6.084 0.756 ; 
        RECT 5.472 0.252 6.084 0.324 ; 
        RECT 5.472 0.252 5.544 0.756 ; 
        RECT 4.392 0.252 4.464 0.756 ; 
        RECT 4.244 0.252 4.464 0.324 ; 
        RECT 3.744 0.252 3.964 0.324 ; 
        RECT 3.744 0.252 3.816 0.756 ; 
        RECT 2.664 0.252 2.736 0.756 ; 
        RECT 2.512 0.252 2.736 0.324 ; 
        RECT 2.016 0.252 2.236 0.324 ; 
        RECT 2.016 0.252 2.088 0.756 ; 
        RECT 0.936 0.252 1.008 0.756 ; 
        RECT 0.784 0.252 1.008 0.324 ; 
        RECT 0.228 0.108 0.488 0.18 ; 
        RECT 0.228 0.108 0.3 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 5.04 0.396 5.264 0.468 ; 
      RECT 5.04 0.252 5.112 0.468 ; 
      RECT 4.696 0.252 5.304 0.324 ; 
      RECT 4.62 0.54 5.24 0.612 ; 
      RECT 4.824 0.396 4.896 0.612 ; 
      RECT 4.664 0.396 4.896 0.468 ; 
      RECT 2.968 0.54 3.588 0.612 ; 
      RECT 3.312 0.396 3.384 0.612 ; 
      RECT 3.312 0.396 3.544 0.468 ; 
      RECT 2.944 0.396 3.168 0.468 ; 
      RECT 3.096 0.252 3.168 0.468 ; 
      RECT 2.904 0.252 3.512 0.324 ; 
      RECT 1.24 0.54 1.86 0.612 ; 
      RECT 1.584 0.396 1.656 0.612 ; 
      RECT 1.584 0.396 1.816 0.468 ; 
      RECT 1.216 0.396 1.44 0.468 ; 
      RECT 1.368 0.252 1.44 0.468 ; 
      RECT 1.176 0.252 1.784 0.324 ; 
  END 
END CKINVDCx16_ASAP7_6t_SL 


MACRO CKINVDCx20_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN CKINVDCx20_ASAP7_6t_SL 0 0 ; 
  SIZE 8.208 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 7.372 0.396 7.748 0.468 ; 
        RECT 7.52 0.108 7.616 0.468 ; 
        RECT 0.592 0.108 7.616 0.18 ; 
        RECT 5.648 0.396 6.02 0.468 ; 
        RECT 5.796 0.108 5.868 0.468 ; 
        RECT 3.92 0.396 4.288 0.468 ; 
        RECT 4.068 0.108 4.14 0.468 ; 
        RECT 2.188 0.396 2.56 0.468 ; 
        RECT 2.34 0.108 2.412 0.468 ; 
        RECT 0.504 0.396 0.832 0.468 ; 
        RECT 0.592 0.108 0.684 0.468 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 8.208 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 8.208 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.16 0.684 8.048 0.756 ; 
        RECT 7.976 0.108 8.048 0.756 ; 
        RECT 7.72 0.108 8.048 0.18 ; 
        RECT 7.2 0.252 7.42 0.324 ; 
        RECT 7.2 0.252 7.272 0.756 ; 
        RECT 6.12 0.252 6.192 0.756 ; 
        RECT 5.972 0.252 6.192 0.324 ; 
        RECT 5.472 0.252 5.692 0.324 ; 
        RECT 5.472 0.252 5.544 0.756 ; 
        RECT 4.392 0.252 4.464 0.756 ; 
        RECT 4.244 0.252 4.464 0.324 ; 
        RECT 3.744 0.252 3.964 0.324 ; 
        RECT 3.744 0.252 3.816 0.756 ; 
        RECT 2.664 0.252 2.736 0.756 ; 
        RECT 2.516 0.252 2.736 0.324 ; 
        RECT 2.016 0.252 2.236 0.324 ; 
        RECT 2.016 0.252 2.088 0.756 ; 
        RECT 0.936 0.252 1.008 0.756 ; 
        RECT 0.788 0.252 1.008 0.324 ; 
        RECT 0.16 0.108 0.488 0.18 ; 
        RECT 0.16 0.108 0.232 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 6.768 0.396 6.992 0.468 ; 
      RECT 6.768 0.252 6.84 0.468 ; 
      RECT 6.424 0.252 7.032 0.324 ; 
      RECT 6.348 0.54 6.968 0.612 ; 
      RECT 6.552 0.396 6.624 0.612 ; 
      RECT 6.392 0.396 6.624 0.468 ; 
      RECT 5.04 0.396 5.264 0.468 ; 
      RECT 5.04 0.252 5.112 0.468 ; 
      RECT 4.696 0.252 5.304 0.324 ; 
      RECT 4.62 0.54 5.24 0.612 ; 
      RECT 4.824 0.396 4.896 0.612 ; 
      RECT 4.664 0.396 4.896 0.468 ; 
      RECT 2.968 0.54 3.588 0.612 ; 
      RECT 3.312 0.396 3.384 0.612 ; 
      RECT 3.312 0.396 3.544 0.468 ; 
      RECT 2.944 0.396 3.168 0.468 ; 
      RECT 3.096 0.252 3.168 0.468 ; 
      RECT 2.904 0.252 3.512 0.324 ; 
      RECT 1.24 0.54 1.86 0.612 ; 
      RECT 1.584 0.396 1.656 0.612 ; 
      RECT 1.584 0.396 1.816 0.468 ; 
      RECT 1.216 0.396 1.44 0.468 ; 
      RECT 1.368 0.252 1.44 0.468 ; 
      RECT 1.176 0.252 1.784 0.324 ; 
  END 
END CKINVDCx20_ASAP7_6t_SL 


MACRO CKINVDCx5p5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN CKINVDCx5p5_ASAP7_6t_SL 0 0 ; 
  SIZE 4.536 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.048 0.396 4.336 0.468 ; 
        RECT 4.264 0.108 4.336 0.468 ; 
        RECT 0.376 0.108 4.336 0.18 ; 
        RECT 2.752 0.396 3.04 0.468 ; 
        RECT 2.968 0.108 3.04 0.468 ; 
        RECT 1.28 0.396 1.568 0.468 ; 
        RECT 1.28 0.108 1.352 0.468 ; 
        RECT 0.268 0.396 0.448 0.468 ; 
        RECT 0.376 0.108 0.448 0.468 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 4.536 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.536 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.092 0.684 4.16 0.756 ; 
        RECT 3.876 0.252 4.16 0.324 ; 
        RECT 3.876 0.252 3.948 0.756 ; 
        RECT 2.58 0.252 2.864 0.324 ; 
        RECT 2.58 0.252 2.652 0.756 ; 
        RECT 1.668 0.252 1.74 0.756 ; 
        RECT 1.456 0.252 1.74 0.324 ; 
        RECT 0.092 0.108 0.272 0.18 ; 
        RECT 0.092 0.108 0.168 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 3.528 0.396 3.752 0.468 ; 
      RECT 3.528 0.252 3.6 0.468 ; 
      RECT 3.184 0.252 3.776 0.324 ; 
      RECT 3.108 0.54 3.728 0.612 ; 
      RECT 3.312 0.396 3.384 0.612 ; 
      RECT 3.152 0.396 3.384 0.468 ; 
      RECT 1.888 0.54 2.464 0.612 ; 
      RECT 2.232 0.396 2.304 0.612 ; 
      RECT 2.232 0.396 2.464 0.468 ; 
      RECT 1.864 0.396 2.088 0.468 ; 
      RECT 2.016 0.252 2.088 0.468 ; 
      RECT 1.852 0.252 2.432 0.324 ; 
      RECT 0.592 0.54 1.212 0.612 ; 
      RECT 0.936 0.396 1.008 0.612 ; 
      RECT 0.936 0.396 1.168 0.468 ; 
      RECT 0.568 0.396 0.792 0.468 ; 
      RECT 0.72 0.252 0.792 0.468 ; 
      RECT 0.568 0.252 1.136 0.324 ; 
  END 
END CKINVDCx5p5_ASAP7_6t_SL 


MACRO CKINVDCx6p5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN CKINVDCx6p5_ASAP7_6t_SL 0 0 ; 
  SIZE 4.968 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.284 0.396 4.652 0.468 ; 
        RECT 0.16 0.108 4.592 0.18 ; 
        RECT 4.48 0.108 4.552 0.468 ; 
        RECT 2.988 0.396 3.256 0.468 ; 
        RECT 3.184 0.108 3.256 0.468 ; 
        RECT 1.496 0.396 1.764 0.468 ; 
        RECT 1.496 0.108 1.568 0.468 ; 
        RECT 0.16 0.396 0.468 0.468 ; 
        RECT 0.16 0.108 0.272 0.468 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 4.968 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.968 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 4.864 0.756 ; 
        RECT 4.792 0.252 4.864 0.756 ; 
        RECT 4.696 0.252 4.864 0.324 ; 
        RECT 4.112 0.252 4.376 0.324 ; 
        RECT 4.112 0.252 4.184 0.756 ; 
        RECT 2.808 0.252 3.08 0.324 ; 
        RECT 2.808 0.252 2.88 0.756 ; 
        RECT 1.868 0.252 1.94 0.756 ; 
        RECT 1.672 0.252 1.94 0.324 ; 
        RECT 0.576 0.252 0.648 0.756 ; 
        RECT 0.376 0.252 0.648 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 3.744 0.396 3.968 0.468 ; 
      RECT 3.744 0.252 3.816 0.468 ; 
      RECT 3.4 0.252 4.008 0.324 ; 
      RECT 3.324 0.54 3.944 0.612 ; 
      RECT 3.528 0.396 3.6 0.612 ; 
      RECT 3.368 0.396 3.6 0.468 ; 
      RECT 2.104 0.54 2.704 0.612 ; 
      RECT 2.448 0.396 2.52 0.612 ; 
      RECT 2.448 0.396 2.68 0.468 ; 
      RECT 2.08 0.396 2.304 0.468 ; 
      RECT 2.232 0.252 2.304 0.468 ; 
      RECT 2.044 0.252 2.648 0.324 ; 
      RECT 0.808 0.54 1.428 0.612 ; 
      RECT 1.152 0.396 1.224 0.612 ; 
      RECT 1.152 0.396 1.384 0.468 ; 
      RECT 0.784 0.396 1.008 0.468 ; 
      RECT 0.936 0.252 1.008 0.468 ; 
      RECT 0.756 0.252 1.352 0.324 ; 
  END 
END CKINVDCx6p5_ASAP7_6t_SL 


MACRO CKINVDCx8_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN CKINVDCx8_ASAP7_6t_SL 0 0 ; 
  SIZE 4.752 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.072 0.396 4.36 0.468 ; 
        RECT 4.072 0.108 4.144 0.468 ; 
        RECT 0.108 0.108 4.144 0.18 ; 
        RECT 2.988 0.396 3.268 0.468 ; 
        RECT 3.196 0.108 3.268 0.468 ; 
        RECT 1.484 0.396 1.764 0.468 ; 
        RECT 1.484 0.108 1.556 0.468 ; 
        RECT 0.108 0.396 0.34 0.468 ; 
        RECT 0.108 0.684 0.272 0.756 ; 
        RECT 0.108 0.108 0.18 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 4.752 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.752 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.684 4.548 0.756 ; 
        RECT 4.476 0.108 4.548 0.756 ; 
        RECT 4.264 0.108 4.548 0.18 ; 
        RECT 2.816 0.252 3.084 0.324 ; 
        RECT 2.816 0.252 2.888 0.756 ; 
        RECT 1.864 0.252 1.936 0.756 ; 
        RECT 1.668 0.252 1.936 0.324 ; 
        RECT 0.504 0.252 0.576 0.756 ; 
        RECT 0.376 0.252 0.576 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 3.744 0.396 3.968 0.468 ; 
      RECT 3.744 0.252 3.816 0.468 ; 
      RECT 3.4 0.252 3.972 0.324 ; 
      RECT 3.36 0.54 3.944 0.612 ; 
      RECT 3.528 0.396 3.6 0.612 ; 
      RECT 3.368 0.396 3.6 0.468 ; 
      RECT 2.104 0.54 2.716 0.612 ; 
      RECT 2.448 0.396 2.52 0.612 ; 
      RECT 2.448 0.396 2.68 0.468 ; 
      RECT 2.08 0.396 2.304 0.468 ; 
      RECT 2.232 0.252 2.304 0.468 ; 
      RECT 2.04 0.252 2.648 0.324 ; 
      RECT 0.808 0.54 1.408 0.612 ; 
      RECT 1.152 0.396 1.224 0.612 ; 
      RECT 1.152 0.396 1.384 0.468 ; 
      RECT 0.784 0.396 1.008 0.468 ; 
      RECT 0.936 0.252 1.008 0.468 ; 
      RECT 0.744 0.252 1.352 0.324 ; 
  END 
END CKINVDCx8_ASAP7_6t_SL 


MACRO CKINVDCx9p5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN CKINVDCx9p5_ASAP7_6t_SL 0 0 ; 
  SIZE 6.048 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.148 0.396 5.652 0.468 ; 
        RECT 5.356 0.108 5.456 0.468 ; 
        RECT 0.16 0.108 5.456 0.18 ; 
        RECT 3.42 0.396 3.924 0.468 ; 
        RECT 3.636 0.108 3.708 0.468 ; 
        RECT 1.692 0.396 2.196 0.468 ; 
        RECT 1.904 0.108 1.976 0.468 ; 
        RECT 0.16 0.396 0.468 0.468 ; 
        RECT 0.16 0.108 0.256 0.468 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 6.048 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 6.048 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.16 0.684 5.888 0.756 ; 
        RECT 5.816 0.252 5.888 0.756 ; 
        RECT 5.56 0.252 5.888 0.324 ; 
        RECT 4.976 0.252 5.24 0.324 ; 
        RECT 4.976 0.252 5.048 0.756 ; 
        RECT 4.024 0.252 4.096 0.756 ; 
        RECT 3.832 0.252 4.096 0.324 ; 
        RECT 3.248 0.252 3.512 0.324 ; 
        RECT 3.248 0.252 3.32 0.756 ; 
        RECT 2.296 0.252 2.368 0.756 ; 
        RECT 2.104 0.252 2.368 0.324 ; 
        RECT 1.52 0.252 1.784 0.324 ; 
        RECT 1.52 0.252 1.592 0.756 ; 
        RECT 0.568 0.252 0.64 0.756 ; 
        RECT 0.356 0.252 0.64 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 4.608 0.396 4.832 0.468 ; 
      RECT 4.608 0.252 4.68 0.468 ; 
      RECT 4.264 0.252 4.872 0.324 ; 
      RECT 4.22 0.54 4.808 0.612 ; 
      RECT 4.392 0.396 4.464 0.612 ; 
      RECT 4.232 0.396 4.464 0.468 ; 
      RECT 2.536 0.54 3.12 0.612 ; 
      RECT 2.88 0.396 2.952 0.612 ; 
      RECT 2.88 0.396 3.112 0.468 ; 
      RECT 2.512 0.396 2.736 0.468 ; 
      RECT 2.664 0.252 2.736 0.468 ; 
      RECT 2.472 0.252 3.08 0.324 ; 
      RECT 0.808 0.54 1.392 0.612 ; 
      RECT 1.152 0.396 1.224 0.612 ; 
      RECT 1.152 0.396 1.384 0.468 ; 
      RECT 0.784 0.396 1.008 0.468 ; 
      RECT 0.936 0.252 1.008 0.468 ; 
      RECT 0.744 0.252 1.352 0.324 ; 
  END 
END CKINVDCx9p5_ASAP7_6t_SL 


MACRO DECAPx10_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DECAPx10_ASAP7_6t_SL 0 0 ; 
  SIZE 4.752 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 4.752 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.752 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.232 0.18 2.304 0.468 ; 
      RECT 2.232 0.18 4.592 0.252 ; 
      RECT 0.16 0.612 2.52 0.684 ; 
      RECT 2.448 0.396 2.52 0.684 ; 
  END 
END DECAPx10_ASAP7_6t_SL 


MACRO DECAPx1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DECAPx1_ASAP7_6t_SL 0 0 ; 
  SIZE 0.864 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 0.864 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.864 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.612 0.576 0.684 ; 
      RECT 0.504 0.396 0.576 0.684 ; 
      RECT 0.288 0.18 0.36 0.468 ; 
      RECT 0.288 0.18 0.468 0.252 ; 
  END 
END DECAPx1_ASAP7_6t_SL 


MACRO DECAPx2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DECAPx2_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 0.504 0.18 0.576 0.468 ; 
      RECT 0.504 0.18 1.136 0.252 ; 
      RECT 0.16 0.612 0.792 0.684 ; 
      RECT 0.72 0.396 0.792 0.684 ; 
  END 
END DECAPx2_ASAP7_6t_SL 


MACRO DECAPx2b_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DECAPx2b_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.54 0.996 0.612 ; 
      RECT 0.72 0.396 0.792 0.612 ; 
      RECT 0.72 0.396 0.952 0.468 ; 
      RECT 0.352 0.396 0.576 0.468 ; 
      RECT 0.504 0.252 0.576 0.468 ; 
      RECT 0.312 0.252 0.92 0.324 ; 
  END 
END DECAPx2b_ASAP7_6t_SL 


MACRO DECAPx4_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DECAPx4_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 0.936 0.18 1.008 0.468 ; 
      RECT 0.936 0.18 2 0.252 ; 
      RECT 0.16 0.612 1.224 0.684 ; 
      RECT 1.152 0.396 1.224 0.684 ; 
  END 
END DECAPx4_ASAP7_6t_SL 


MACRO DECAPx6_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DECAPx6_ASAP7_6t_SL 0 0 ; 
  SIZE 3.024 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.024 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.024 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 1.368 0.18 1.44 0.468 ; 
      RECT 1.368 0.18 2.864 0.252 ; 
      RECT 0.16 0.612 1.656 0.684 ; 
      RECT 1.584 0.396 1.656 0.684 ; 
  END 
END DECAPx6_ASAP7_6t_SL 


MACRO DFFARHQNx1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFFARHQNx1_ASAP7_6t_SL 0 0 ; 
  SIZE 5.184 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.208 0.684 0.54 0.756 ; 
        RECT 0.208 0.108 0.54 0.18 ; 
        RECT 0.208 0.396 0.36 0.468 ; 
        RECT 0.208 0.108 0.28 0.756 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.08 0.108 1.38 0.18 ; 
        RECT 0.764 0.684 1.236 0.756 ; 
        RECT 1.08 0.396 1.224 0.468 ; 
        RECT 1.08 0.108 1.152 0.756 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.852 0.684 5.112 0.756 ; 
        RECT 5.04 0.108 5.112 0.756 ; 
        RECT 4.852 0.108 5.112 0.18 ; 
    END 
  END QN 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 5.184 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.184 0.036 ; 
    END 
  END VSS 
  PIN RESETN 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 2.104 0.108 4.592 0.18 ; 
      LAYER M1 ; 
        RECT 4.444 0.108 4.608 0.18 ; 
        RECT 4.444 0.108 4.516 0.392 ; 
        RECT 2.02 0.108 2.244 0.18 ; 
        RECT 2.02 0.108 2.092 0.352 ; 
      LAYER V1 ; 
        RECT 2.124 0.108 2.196 0.18 ; 
        RECT 4.5 0.108 4.572 0.18 ; 
    END 
  END RESETN 
  OBS 
    LAYER M1 ; 
      RECT 4.824 0.252 4.896 0.5 ; 
      RECT 4.768 0.252 4.916 0.324 ; 
      RECT 4.276 0.684 4.596 0.756 ; 
      RECT 4.276 0.108 4.348 0.756 ; 
      RECT 3.744 0.108 3.816 0.352 ; 
      RECT 3.744 0.108 4.348 0.18 ; 
      RECT 3.816 0.54 3.952 0.612 ; 
      RECT 3.816 0.452 3.896 0.612 ; 
      RECT 3.628 0.452 3.896 0.524 ; 
      RECT 3.42 0.52 3.492 0.7 ; 
      RECT 3.456 0.108 3.528 0.604 ; 
      RECT 3.456 0.252 3.616 0.324 ; 
      RECT 3.184 0.108 3.528 0.18 ; 
      RECT 3.312 0.252 3.384 0.416 ; 
      RECT 3.232 0.252 3.384 0.324 ; 
      RECT 2.996 0.684 3.296 0.756 ; 
      RECT 2.996 0.108 3.068 0.756 ; 
      RECT 2.456 0.108 2.528 0.528 ; 
      RECT 2.456 0.108 3.068 0.18 ; 
      RECT 3.14 0.54 3.288 0.612 ; 
      RECT 3.14 0.432 3.212 0.612 ; 
      RECT 2.168 0.54 2.32 0.612 ; 
      RECT 2.012 0.476 2.276 0.548 ; 
      RECT 1.416 0.684 1.796 0.756 ; 
      RECT 1.724 0.216 1.796 0.756 ; 
      RECT 1.572 0.252 1.644 0.504 ; 
      RECT 1.496 0.252 1.644 0.324 ; 
      RECT 1.288 0.54 1.44 0.612 ; 
      RECT 1.368 0.392 1.44 0.612 ; 
      RECT 0.728 0.54 1.008 0.612 ; 
      RECT 0.936 0.252 1.008 0.612 ; 
      RECT 0.78 0.252 1.008 0.324 ; 
      RECT 0.504 0.252 0.576 0.504 ; 
      RECT 0.444 0.252 0.616 0.324 ; 
      RECT 2.64 0.396 2.876 0.468 ; 
      RECT 1.908 0.684 2.492 0.756 ; 
      RECT 0.064 0.196 0.136 0.668 ; 
    LAYER M2 ; 
      RECT 3.528 0.252 4.916 0.324 ; 
      RECT 0.808 0.54 3.944 0.612 ; 
      RECT 0.064 0.252 3.356 0.324 ; 
      RECT 1.704 0.396 2.816 0.468 ; 
    LAYER V1 ; 
      RECT 4.824 0.252 4.896 0.324 ; 
      RECT 3.852 0.54 3.924 0.612 ; 
      RECT 3.528 0.252 3.6 0.324 ; 
      RECT 3.284 0.252 3.356 0.324 ; 
      RECT 3.16 0.54 3.232 0.612 ; 
      RECT 2.704 0.396 2.776 0.468 ; 
      RECT 2.204 0.54 2.276 0.612 ; 
      RECT 1.724 0.396 1.796 0.468 ; 
      RECT 1.54 0.252 1.612 0.324 ; 
      RECT 1.332 0.54 1.404 0.612 ; 
      RECT 0.828 0.54 0.9 0.612 ; 
      RECT 0.504 0.252 0.576 0.324 ; 
      RECT 0.064 0.252 0.136 0.324 ; 
  END 
END DFFARHQNx1_ASAP7_6t_SL 


MACRO DFFASHQNx1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFFASHQNx1_ASAP7_6t_SL 0 0 ; 
  SIZE 5.184 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.208 0.684 0.54 0.756 ; 
        RECT 0.208 0.108 0.54 0.18 ; 
        RECT 0.208 0.396 0.36 0.468 ; 
        RECT 0.208 0.108 0.28 0.756 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.08 0.108 1.38 0.18 ; 
        RECT 0.764 0.684 1.236 0.756 ; 
        RECT 1.08 0.396 1.224 0.468 ; 
        RECT 1.08 0.108 1.152 0.756 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.852 0.684 5.112 0.756 ; 
        RECT 5.04 0.108 5.112 0.756 ; 
        RECT 4.852 0.108 5.112 0.18 ; 
    END 
  END QN 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 5.184 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.184 0.036 ; 
    END 
  END VSS 
  PIN SETN 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 2.832 0.396 4.368 0.468 ; 
      LAYER M1 ; 
        RECT 4.276 0.28 4.348 0.568 ; 
        RECT 3.96 0.28 4.348 0.352 ; 
        RECT 2.736 0.684 2.924 0.756 ; 
        RECT 2.852 0.376 2.924 0.756 ; 
      LAYER V1 ; 
        RECT 2.852 0.396 2.924 0.468 ; 
        RECT 4.276 0.396 4.348 0.468 ; 
    END 
  END SETN 
  OBS 
    LAYER M1 ; 
      RECT 4.824 0.252 4.896 0.5 ; 
      RECT 4.768 0.252 4.916 0.324 ; 
      RECT 4.264 0.684 4.56 0.756 ; 
      RECT 4.488 0.108 4.56 0.756 ; 
      RECT 3.744 0.108 3.816 0.352 ; 
      RECT 3.744 0.108 4.56 0.18 ; 
      RECT 3.816 0.54 4.088 0.612 ; 
      RECT 3.816 0.452 3.896 0.612 ; 
      RECT 3.628 0.452 3.896 0.524 ; 
      RECT 3.42 0.52 3.492 0.7 ; 
      RECT 3.456 0.108 3.528 0.604 ; 
      RECT 3.456 0.252 3.616 0.324 ; 
      RECT 3.184 0.108 3.528 0.18 ; 
      RECT 3.312 0.252 3.384 0.416 ; 
      RECT 3.232 0.252 3.384 0.324 ; 
      RECT 2.996 0.684 3.296 0.756 ; 
      RECT 2.996 0.108 3.068 0.756 ; 
      RECT 2.24 0.54 2.648 0.612 ; 
      RECT 2.24 0.108 2.312 0.612 ; 
      RECT 2.24 0.108 3.068 0.18 ; 
      RECT 3.14 0.54 3.288 0.612 ; 
      RECT 3.14 0.432 3.212 0.612 ; 
      RECT 1.868 0.54 2.104 0.612 ; 
      RECT 1.868 0.432 1.94 0.612 ; 
      RECT 1.416 0.684 1.796 0.756 ; 
      RECT 1.724 0.216 1.796 0.756 ; 
      RECT 1.572 0.252 1.644 0.504 ; 
      RECT 1.496 0.252 1.644 0.324 ; 
      RECT 1.288 0.54 1.44 0.612 ; 
      RECT 1.368 0.392 1.44 0.612 ; 
      RECT 0.728 0.54 1.008 0.612 ; 
      RECT 0.936 0.252 1.008 0.612 ; 
      RECT 0.78 0.252 1.008 0.324 ; 
      RECT 0.504 0.252 0.576 0.504 ; 
      RECT 0.444 0.252 0.616 0.324 ; 
      RECT 3.616 0.684 4.14 0.756 ; 
      RECT 2.424 0.396 2.66 0.468 ; 
      RECT 0.064 0.196 0.136 0.668 ; 
    LAYER M2 ; 
      RECT 3.528 0.252 4.924 0.324 ; 
      RECT 0.808 0.54 4.052 0.612 ; 
      RECT 0.064 0.252 3.356 0.324 ; 
      RECT 1.704 0.396 2.6 0.468 ; 
    LAYER V1 ; 
      RECT 4.824 0.252 4.896 0.324 ; 
      RECT 3.96 0.54 4.032 0.612 ; 
      RECT 3.528 0.252 3.6 0.324 ; 
      RECT 3.284 0.252 3.356 0.324 ; 
      RECT 3.16 0.54 3.232 0.612 ; 
      RECT 2.488 0.396 2.56 0.468 ; 
      RECT 1.988 0.54 2.06 0.612 ; 
      RECT 1.724 0.396 1.796 0.468 ; 
      RECT 1.54 0.252 1.612 0.324 ; 
      RECT 1.332 0.54 1.404 0.612 ; 
      RECT 0.828 0.54 0.9 0.612 ; 
      RECT 0.504 0.252 0.576 0.324 ; 
      RECT 0.064 0.252 0.136 0.324 ; 
  END 
END DFFASHQNx1_ASAP7_6t_SL 


MACRO DFFASRHQNx1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFFASRHQNx1_ASAP7_6t_SL 0 0 ; 
  SIZE 5.616 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.208 0.684 0.54 0.756 ; 
        RECT 0.208 0.108 0.54 0.18 ; 
        RECT 0.208 0.396 0.36 0.468 ; 
        RECT 0.208 0.108 0.28 0.756 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.08 0.108 1.38 0.18 ; 
        RECT 0.764 0.684 1.236 0.756 ; 
        RECT 1.08 0.396 1.224 0.468 ; 
        RECT 1.08 0.108 1.152 0.756 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.284 0.684 5.544 0.756 ; 
        RECT 5.472 0.108 5.544 0.756 ; 
        RECT 5.284 0.108 5.544 0.18 ; 
    END 
  END QN 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 5.616 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.616 0.036 ; 
    END 
  END VSS 
  PIN RESETN 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 2.104 0.108 5.024 0.18 ; 
      LAYER M1 ; 
        RECT 4.876 0.108 5.04 0.18 ; 
        RECT 4.876 0.108 4.948 0.392 ; 
        RECT 2.02 0.108 2.244 0.18 ; 
        RECT 2.02 0.108 2.092 0.352 ; 
      LAYER V1 ; 
        RECT 2.124 0.108 2.196 0.18 ; 
        RECT 4.932 0.108 5.004 0.18 ; 
    END 
  END RESETN 
  PIN SETN 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 3.048 0.396 4.656 0.468 ; 
      LAYER M1 ; 
        RECT 4.564 0.28 4.636 0.568 ; 
        RECT 4.176 0.28 4.636 0.352 ; 
        RECT 2.952 0.684 3.14 0.756 ; 
        RECT 3.068 0.376 3.14 0.756 ; 
      LAYER V1 ; 
        RECT 3.068 0.396 3.14 0.468 ; 
        RECT 4.564 0.396 4.636 0.468 ; 
    END 
  END SETN 
  OBS 
    LAYER M1 ; 
      RECT 5.256 0.252 5.328 0.5 ; 
      RECT 5.2 0.252 5.348 0.324 ; 
      RECT 4.708 0.684 5.028 0.756 ; 
      RECT 4.708 0.108 4.78 0.756 ; 
      RECT 3.96 0.108 4.032 0.352 ; 
      RECT 3.96 0.108 4.78 0.18 ; 
      RECT 4.032 0.54 4.304 0.612 ; 
      RECT 4.032 0.452 4.112 0.612 ; 
      RECT 3.844 0.452 4.112 0.524 ; 
      RECT 3.636 0.52 3.708 0.7 ; 
      RECT 3.672 0.108 3.744 0.604 ; 
      RECT 3.672 0.252 3.832 0.324 ; 
      RECT 3.4 0.108 3.744 0.18 ; 
      RECT 3.528 0.252 3.6 0.416 ; 
      RECT 3.448 0.252 3.6 0.324 ; 
      RECT 3.212 0.684 3.512 0.756 ; 
      RECT 3.212 0.108 3.284 0.756 ; 
      RECT 2.456 0.54 2.864 0.612 ; 
      RECT 2.456 0.108 2.528 0.612 ; 
      RECT 2.456 0.108 3.284 0.18 ; 
      RECT 3.356 0.54 3.504 0.612 ; 
      RECT 3.356 0.432 3.428 0.612 ; 
      RECT 2.168 0.54 2.32 0.612 ; 
      RECT 2.012 0.476 2.276 0.548 ; 
      RECT 1.416 0.684 1.796 0.756 ; 
      RECT 1.724 0.216 1.796 0.756 ; 
      RECT 1.572 0.252 1.644 0.504 ; 
      RECT 1.496 0.252 1.644 0.324 ; 
      RECT 1.288 0.54 1.44 0.612 ; 
      RECT 1.368 0.392 1.44 0.612 ; 
      RECT 0.728 0.54 1.008 0.612 ; 
      RECT 0.936 0.252 1.008 0.612 ; 
      RECT 0.78 0.252 1.008 0.324 ; 
      RECT 0.504 0.252 0.576 0.504 ; 
      RECT 0.444 0.252 0.616 0.324 ; 
      RECT 3.832 0.684 4.376 0.756 ; 
      RECT 2.64 0.396 2.876 0.468 ; 
      RECT 1.908 0.684 2.492 0.756 ; 
      RECT 0.064 0.196 0.136 0.668 ; 
    LAYER M2 ; 
      RECT 3.744 0.252 5.348 0.324 ; 
      RECT 0.808 0.54 4.268 0.612 ; 
      RECT 0.064 0.252 3.572 0.324 ; 
      RECT 1.704 0.396 2.816 0.468 ; 
    LAYER V1 ; 
      RECT 5.256 0.252 5.328 0.324 ; 
      RECT 4.176 0.54 4.248 0.612 ; 
      RECT 3.744 0.252 3.816 0.324 ; 
      RECT 3.5 0.252 3.572 0.324 ; 
      RECT 3.376 0.54 3.448 0.612 ; 
      RECT 2.704 0.396 2.776 0.468 ; 
      RECT 2.204 0.54 2.276 0.612 ; 
      RECT 1.724 0.396 1.796 0.468 ; 
      RECT 1.54 0.252 1.612 0.324 ; 
      RECT 1.332 0.54 1.404 0.612 ; 
      RECT 0.828 0.54 0.9 0.612 ; 
      RECT 0.504 0.252 0.576 0.324 ; 
      RECT 0.064 0.252 0.136 0.324 ; 
  END 
END DFFASRHQNx1_ASAP7_6t_SL 


MACRO DFFHQNx1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFFHQNx1_ASAP7_6t_SL 0 0 ; 
  SIZE 4.32 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.704 0.756 ; 
        RECT 0.376 0.108 0.704 0.18 ; 
        RECT 0.376 0.512 0.468 0.756 ; 
        RECT 0.288 0.26 0.46 0.332 ; 
        RECT 0.376 0.108 0.46 0.332 ; 
        RECT 0.288 0.512 0.468 0.584 ; 
        RECT 0.288 0.26 0.36 0.584 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.08 0.108 1.568 0.18 ; 
        RECT 1.004 0.684 1.352 0.756 ; 
        RECT 1.08 0.108 1.152 0.756 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 3.812 0.684 4.248 0.756 ; 
        RECT 4.176 0.108 4.248 0.756 ; 
        RECT 3.812 0.108 4.248 0.18 ; 
    END 
  END QN 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 4.32 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.32 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 3.524 0.252 3.596 0.504 ; 
      RECT 3.448 0.252 3.596 0.324 ; 
      RECT 3.24 0.684 3.512 0.756 ; 
      RECT 3.24 0.108 3.312 0.756 ; 
      RECT 3.076 0.28 3.312 0.352 ; 
      RECT 3.236 0.108 3.312 0.352 ; 
      RECT 3.236 0.108 3.512 0.18 ; 
      RECT 2.752 0.68 2.952 0.752 ; 
      RECT 2.88 0.108 2.952 0.752 ; 
      RECT 2.536 0.108 2.952 0.18 ; 
      RECT 2.664 0.252 2.736 0.492 ; 
      RECT 2.616 0.252 2.776 0.324 ; 
      RECT 2.404 0.54 2.56 0.612 ; 
      RECT 2.448 0.376 2.52 0.612 ; 
      RECT 2.088 0.684 2.512 0.756 ; 
      RECT 2.088 0.188 2.16 0.756 ; 
      RECT 1.976 0.308 2.16 0.38 ; 
      RECT 2.088 0.188 2.412 0.26 ; 
      RECT 1.476 0.684 1.856 0.756 ; 
      RECT 1.784 0.108 1.856 0.756 ; 
      RECT 1.692 0.108 1.856 0.18 ; 
      RECT 1.584 0.252 1.656 0.504 ; 
      RECT 1.508 0.252 1.656 0.324 ; 
      RECT 1.224 0.54 1.508 0.612 ; 
      RECT 1.224 0.396 1.296 0.612 ; 
      RECT 1.224 0.396 1.472 0.468 ; 
      RECT 0.804 0.448 0.876 0.632 ; 
      RECT 0.804 0.448 0.976 0.52 ; 
      RECT 0.9 0.108 0.976 0.52 ; 
      RECT 0.828 0.108 0.976 0.18 ; 
      RECT 0.572 0.252 0.644 0.468 ; 
      RECT 0.572 0.252 0.732 0.324 ; 
      RECT 0.064 0.684 0.272 0.756 ; 
      RECT 0.064 0.108 0.136 0.756 ; 
      RECT 0.064 0.108 0.252 0.18 ; 
      RECT 3.096 0.452 3.168 0.688 ; 
      RECT 2.232 0.376 2.304 0.576 ; 
      RECT 1.944 0.504 2.016 0.688 ; 
    LAYER M2 ; 
      RECT 2.88 0.252 3.596 0.324 ; 
      RECT 0.784 0.54 3.188 0.612 ; 
      RECT 0.064 0.252 2.736 0.324 ; 
      RECT 1.784 0.396 2.304 0.468 ; 
    LAYER V1 ; 
      RECT 3.504 0.252 3.576 0.324 ; 
      RECT 3.096 0.54 3.168 0.612 ; 
      RECT 2.88 0.252 2.952 0.324 ; 
      RECT 2.664 0.252 2.736 0.324 ; 
      RECT 2.448 0.54 2.52 0.612 ; 
      RECT 2.232 0.396 2.304 0.468 ; 
      RECT 1.944 0.54 2.016 0.612 ; 
      RECT 1.784 0.396 1.856 0.468 ; 
      RECT 1.564 0.252 1.636 0.324 ; 
      RECT 1.26 0.54 1.332 0.612 ; 
      RECT 0.804 0.54 0.876 0.612 ; 
      RECT 0.612 0.252 0.684 0.324 ; 
      RECT 0.064 0.252 0.136 0.324 ; 
  END 
END DFFHQNx1_ASAP7_6t_SL 


MACRO DFFHQNx2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFFHQNx2_ASAP7_6t_SL 0 0 ; 
  SIZE 4.536 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.704 0.756 ; 
        RECT 0.376 0.108 0.704 0.18 ; 
        RECT 0.376 0.512 0.468 0.756 ; 
        RECT 0.288 0.26 0.46 0.332 ; 
        RECT 0.376 0.108 0.46 0.332 ; 
        RECT 0.288 0.512 0.468 0.584 ; 
        RECT 0.288 0.26 0.36 0.584 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.08 0.108 1.568 0.18 ; 
        RECT 1.004 0.684 1.352 0.756 ; 
        RECT 1.08 0.108 1.152 0.756 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 3.804 0.684 4.248 0.756 ; 
        RECT 4.176 0.108 4.248 0.756 ; 
        RECT 3.804 0.108 4.248 0.18 ; 
    END 
  END QN 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 4.536 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.536 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 3.524 0.252 3.596 0.504 ; 
      RECT 3.448 0.252 3.596 0.324 ; 
      RECT 3.24 0.684 3.512 0.756 ; 
      RECT 3.24 0.108 3.312 0.756 ; 
      RECT 3.076 0.28 3.312 0.352 ; 
      RECT 3.236 0.108 3.312 0.352 ; 
      RECT 3.236 0.108 3.512 0.18 ; 
      RECT 2.752 0.68 2.952 0.752 ; 
      RECT 2.88 0.108 2.952 0.752 ; 
      RECT 2.536 0.108 2.952 0.18 ; 
      RECT 2.664 0.252 2.736 0.492 ; 
      RECT 2.616 0.252 2.776 0.324 ; 
      RECT 2.404 0.54 2.56 0.612 ; 
      RECT 2.448 0.376 2.52 0.612 ; 
      RECT 2.088 0.684 2.512 0.756 ; 
      RECT 2.088 0.188 2.16 0.756 ; 
      RECT 1.976 0.308 2.16 0.38 ; 
      RECT 2.088 0.188 2.412 0.26 ; 
      RECT 1.476 0.684 1.856 0.756 ; 
      RECT 1.784 0.108 1.856 0.756 ; 
      RECT 1.692 0.108 1.856 0.18 ; 
      RECT 1.584 0.252 1.656 0.504 ; 
      RECT 1.508 0.252 1.656 0.324 ; 
      RECT 1.224 0.54 1.508 0.612 ; 
      RECT 1.224 0.396 1.296 0.612 ; 
      RECT 1.224 0.396 1.472 0.468 ; 
      RECT 0.804 0.448 0.876 0.632 ; 
      RECT 0.804 0.448 0.976 0.52 ; 
      RECT 0.9 0.108 0.976 0.52 ; 
      RECT 0.828 0.108 0.976 0.18 ; 
      RECT 0.572 0.252 0.644 0.468 ; 
      RECT 0.572 0.252 0.732 0.324 ; 
      RECT 0.064 0.684 0.272 0.756 ; 
      RECT 0.064 0.108 0.136 0.756 ; 
      RECT 0.064 0.108 0.252 0.18 ; 
      RECT 3.096 0.452 3.168 0.688 ; 
      RECT 2.232 0.376 2.304 0.576 ; 
      RECT 1.944 0.504 2.016 0.688 ; 
    LAYER M2 ; 
      RECT 2.88 0.252 3.596 0.324 ; 
      RECT 0.784 0.54 3.188 0.612 ; 
      RECT 0.064 0.252 2.736 0.324 ; 
      RECT 1.784 0.396 2.304 0.468 ; 
    LAYER V1 ; 
      RECT 3.504 0.252 3.576 0.324 ; 
      RECT 3.096 0.54 3.168 0.612 ; 
      RECT 2.88 0.252 2.952 0.324 ; 
      RECT 2.664 0.252 2.736 0.324 ; 
      RECT 2.448 0.54 2.52 0.612 ; 
      RECT 2.232 0.396 2.304 0.468 ; 
      RECT 1.944 0.54 2.016 0.612 ; 
      RECT 1.784 0.396 1.856 0.468 ; 
      RECT 1.564 0.252 1.636 0.324 ; 
      RECT 1.26 0.54 1.332 0.612 ; 
      RECT 0.804 0.54 0.876 0.612 ; 
      RECT 0.612 0.252 0.684 0.324 ; 
      RECT 0.064 0.252 0.136 0.324 ; 
  END 
END DFFHQNx2_ASAP7_6t_SL 


MACRO DFFHQNx3_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFFHQNx3_ASAP7_6t_SL 0 0 ; 
  SIZE 4.752 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.704 0.756 ; 
        RECT 0.376 0.108 0.704 0.18 ; 
        RECT 0.376 0.512 0.468 0.756 ; 
        RECT 0.288 0.26 0.46 0.332 ; 
        RECT 0.376 0.108 0.46 0.332 ; 
        RECT 0.288 0.512 0.468 0.584 ; 
        RECT 0.288 0.26 0.36 0.584 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.08 0.108 1.568 0.18 ; 
        RECT 1.004 0.684 1.352 0.756 ; 
        RECT 1.08 0.108 1.152 0.756 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.044 0.684 4.676 0.756 ; 
        RECT 4.604 0.108 4.676 0.756 ; 
        RECT 4.028 0.108 4.676 0.18 ; 
    END 
  END QN 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 4.752 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.752 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 3.524 0.252 3.596 0.504 ; 
      RECT 3.448 0.252 3.596 0.324 ; 
      RECT 3.24 0.684 3.512 0.756 ; 
      RECT 3.24 0.108 3.312 0.756 ; 
      RECT 3.076 0.28 3.312 0.352 ; 
      RECT 3.236 0.108 3.312 0.352 ; 
      RECT 3.236 0.108 3.512 0.18 ; 
      RECT 2.752 0.68 2.952 0.752 ; 
      RECT 2.88 0.108 2.952 0.752 ; 
      RECT 2.536 0.108 2.952 0.18 ; 
      RECT 2.664 0.252 2.736 0.492 ; 
      RECT 2.616 0.252 2.776 0.324 ; 
      RECT 2.404 0.54 2.56 0.612 ; 
      RECT 2.448 0.376 2.52 0.612 ; 
      RECT 2.088 0.684 2.512 0.756 ; 
      RECT 2.088 0.188 2.16 0.756 ; 
      RECT 1.976 0.308 2.16 0.38 ; 
      RECT 2.088 0.188 2.412 0.26 ; 
      RECT 1.476 0.684 1.856 0.756 ; 
      RECT 1.784 0.108 1.856 0.756 ; 
      RECT 1.692 0.108 1.856 0.18 ; 
      RECT 1.584 0.252 1.656 0.504 ; 
      RECT 1.508 0.252 1.656 0.324 ; 
      RECT 1.224 0.54 1.508 0.612 ; 
      RECT 1.224 0.396 1.296 0.612 ; 
      RECT 1.224 0.396 1.472 0.468 ; 
      RECT 0.804 0.448 0.876 0.632 ; 
      RECT 0.804 0.448 0.976 0.52 ; 
      RECT 0.9 0.108 0.976 0.52 ; 
      RECT 0.828 0.108 0.976 0.18 ; 
      RECT 0.572 0.252 0.644 0.468 ; 
      RECT 0.572 0.252 0.732 0.324 ; 
      RECT 0.064 0.684 0.272 0.756 ; 
      RECT 0.064 0.108 0.136 0.756 ; 
      RECT 0.064 0.108 0.252 0.18 ; 
      RECT 3.096 0.452 3.168 0.688 ; 
      RECT 2.232 0.376 2.304 0.576 ; 
      RECT 1.944 0.504 2.016 0.688 ; 
    LAYER M2 ; 
      RECT 2.88 0.252 3.596 0.324 ; 
      RECT 0.784 0.54 3.188 0.612 ; 
      RECT 0.064 0.252 2.736 0.324 ; 
      RECT 1.784 0.396 2.304 0.468 ; 
    LAYER V1 ; 
      RECT 3.504 0.252 3.576 0.324 ; 
      RECT 3.096 0.54 3.168 0.612 ; 
      RECT 2.88 0.252 2.952 0.324 ; 
      RECT 2.664 0.252 2.736 0.324 ; 
      RECT 2.448 0.54 2.52 0.612 ; 
      RECT 2.232 0.396 2.304 0.468 ; 
      RECT 1.944 0.54 2.016 0.612 ; 
      RECT 1.784 0.396 1.856 0.468 ; 
      RECT 1.564 0.252 1.636 0.324 ; 
      RECT 1.26 0.54 1.332 0.612 ; 
      RECT 0.804 0.54 0.876 0.612 ; 
      RECT 0.612 0.252 0.684 0.324 ; 
      RECT 0.064 0.252 0.136 0.324 ; 
  END 
END DFFHQNx3_ASAP7_6t_SL 


MACRO DFFHQx4_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFFHQx4_ASAP7_6t_SL 0 0 ; 
  SIZE 5.4 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.704 0.756 ; 
        RECT 0.376 0.108 0.704 0.18 ; 
        RECT 0.376 0.512 0.468 0.756 ; 
        RECT 0.288 0.26 0.46 0.332 ; 
        RECT 0.376 0.108 0.46 0.332 ; 
        RECT 0.288 0.512 0.468 0.584 ; 
        RECT 0.288 0.26 0.36 0.584 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.08 0.108 1.568 0.18 ; 
        RECT 1.004 0.684 1.352 0.756 ; 
        RECT 1.08 0.108 1.152 0.756 ; 
    END 
  END D 
  PIN Q 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.5 0.684 5.332 0.756 ; 
        RECT 5.252 0.108 5.332 0.756 ; 
        RECT 4.5 0.108 5.332 0.18 ; 
        RECT 4.5 0.588 4.572 0.756 ; 
        RECT 4.5 0.108 4.572 0.276 ; 
    END 
  END Q 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 5.4 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.4 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 4.048 0.684 4.392 0.756 ; 
      RECT 4.32 0.108 4.392 0.756 ; 
      RECT 4.32 0.4 4.7 0.472 ; 
      RECT 4.048 0.108 4.392 0.18 ; 
      RECT 3.524 0.252 3.596 0.504 ; 
      RECT 3.448 0.252 3.596 0.324 ; 
      RECT 3.24 0.684 3.512 0.756 ; 
      RECT 3.24 0.108 3.312 0.756 ; 
      RECT 3.076 0.28 3.312 0.352 ; 
      RECT 3.236 0.108 3.312 0.352 ; 
      RECT 3.236 0.108 3.512 0.18 ; 
      RECT 2.752 0.68 2.952 0.752 ; 
      RECT 2.88 0.108 2.952 0.752 ; 
      RECT 2.536 0.108 2.952 0.18 ; 
      RECT 2.664 0.252 2.736 0.492 ; 
      RECT 2.616 0.252 2.776 0.324 ; 
      RECT 2.404 0.54 2.56 0.612 ; 
      RECT 2.448 0.376 2.52 0.612 ; 
      RECT 2.088 0.684 2.512 0.756 ; 
      RECT 2.088 0.188 2.16 0.756 ; 
      RECT 1.976 0.308 2.16 0.38 ; 
      RECT 2.088 0.188 2.412 0.26 ; 
      RECT 1.476 0.684 1.856 0.756 ; 
      RECT 1.784 0.108 1.856 0.756 ; 
      RECT 1.692 0.108 1.856 0.18 ; 
      RECT 1.584 0.252 1.656 0.504 ; 
      RECT 1.508 0.252 1.656 0.324 ; 
      RECT 1.224 0.54 1.508 0.612 ; 
      RECT 1.224 0.396 1.296 0.612 ; 
      RECT 1.224 0.396 1.472 0.468 ; 
      RECT 0.804 0.448 0.876 0.632 ; 
      RECT 0.804 0.448 0.976 0.52 ; 
      RECT 0.9 0.108 0.976 0.52 ; 
      RECT 0.828 0.108 0.976 0.18 ; 
      RECT 0.572 0.252 0.644 0.468 ; 
      RECT 0.572 0.252 0.732 0.324 ; 
      RECT 0.064 0.684 0.272 0.756 ; 
      RECT 0.064 0.108 0.136 0.756 ; 
      RECT 0.064 0.108 0.252 0.18 ; 
      RECT 3.096 0.452 3.168 0.688 ; 
      RECT 2.232 0.376 2.304 0.576 ; 
      RECT 1.944 0.504 2.016 0.688 ; 
    LAYER M2 ; 
      RECT 2.88 0.252 3.596 0.324 ; 
      RECT 0.784 0.54 3.188 0.612 ; 
      RECT 0.064 0.252 2.736 0.324 ; 
      RECT 1.784 0.396 2.304 0.468 ; 
    LAYER V1 ; 
      RECT 3.504 0.252 3.576 0.324 ; 
      RECT 3.096 0.54 3.168 0.612 ; 
      RECT 2.88 0.252 2.952 0.324 ; 
      RECT 2.664 0.252 2.736 0.324 ; 
      RECT 2.448 0.54 2.52 0.612 ; 
      RECT 2.232 0.396 2.304 0.468 ; 
      RECT 1.944 0.54 2.016 0.612 ; 
      RECT 1.784 0.396 1.856 0.468 ; 
      RECT 1.564 0.252 1.636 0.324 ; 
      RECT 1.26 0.54 1.332 0.612 ; 
      RECT 0.804 0.54 0.876 0.612 ; 
      RECT 0.612 0.252 0.684 0.324 ; 
      RECT 0.064 0.252 0.136 0.324 ; 
  END 
END DFFHQx4_ASAP7_6t_SL 


MACRO DFFLQNx1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFFLQNx1_ASAP7_6t_SL 0 0 ; 
  SIZE 4.32 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.704 0.756 ; 
        RECT 0.376 0.108 0.704 0.18 ; 
        RECT 0.288 0.28 0.468 0.352 ; 
        RECT 0.376 0.108 0.468 0.352 ; 
        RECT 0.376 0.532 0.46 0.756 ; 
        RECT 0.288 0.532 0.46 0.604 ; 
        RECT 0.288 0.28 0.36 0.604 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.08 0.684 1.568 0.756 ; 
        RECT 1.004 0.108 1.352 0.18 ; 
        RECT 1.08 0.108 1.152 0.756 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 3.812 0.684 4.248 0.756 ; 
        RECT 4.176 0.108 4.248 0.756 ; 
        RECT 3.812 0.108 4.248 0.18 ; 
    END 
  END QN 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 4.32 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.32 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 3.448 0.54 3.596 0.612 ; 
      RECT 3.524 0.36 3.596 0.612 ; 
      RECT 3.236 0.684 3.512 0.756 ; 
      RECT 3.236 0.512 3.312 0.756 ; 
      RECT 3.24 0.108 3.312 0.756 ; 
      RECT 3.076 0.512 3.312 0.584 ; 
      RECT 3.24 0.108 3.512 0.18 ; 
      RECT 2.536 0.684 2.952 0.756 ; 
      RECT 2.88 0.112 2.952 0.756 ; 
      RECT 2.752 0.112 2.952 0.184 ; 
      RECT 2.616 0.54 2.776 0.612 ; 
      RECT 2.664 0.372 2.736 0.612 ; 
      RECT 2.448 0.252 2.52 0.488 ; 
      RECT 2.404 0.252 2.56 0.324 ; 
      RECT 2.088 0.604 2.412 0.676 ; 
      RECT 2.088 0.108 2.16 0.676 ; 
      RECT 1.976 0.484 2.16 0.556 ; 
      RECT 2.088 0.108 2.512 0.18 ; 
      RECT 1.692 0.684 1.856 0.756 ; 
      RECT 1.784 0.108 1.856 0.756 ; 
      RECT 1.476 0.108 1.856 0.18 ; 
      RECT 1.508 0.54 1.656 0.612 ; 
      RECT 1.584 0.36 1.656 0.612 ; 
      RECT 1.224 0.396 1.472 0.468 ; 
      RECT 1.224 0.252 1.296 0.468 ; 
      RECT 1.224 0.252 1.508 0.324 ; 
      RECT 0.828 0.684 0.976 0.756 ; 
      RECT 0.9 0.344 0.976 0.756 ; 
      RECT 0.804 0.344 0.976 0.416 ; 
      RECT 0.804 0.232 0.876 0.416 ; 
      RECT 0.572 0.54 0.732 0.612 ; 
      RECT 0.572 0.396 0.644 0.612 ; 
      RECT 0.064 0.684 0.252 0.756 ; 
      RECT 0.064 0.108 0.136 0.756 ; 
      RECT 0.064 0.108 0.272 0.18 ; 
      RECT 3.096 0.176 3.168 0.412 ; 
      RECT 2.232 0.288 2.304 0.488 ; 
      RECT 1.944 0.176 2.016 0.36 ; 
    LAYER M2 ; 
      RECT 2.88 0.54 3.596 0.612 ; 
      RECT 0.784 0.252 3.188 0.324 ; 
      RECT 0.064 0.54 2.736 0.612 ; 
      RECT 1.784 0.396 2.304 0.468 ; 
    LAYER V1 ; 
      RECT 3.504 0.54 3.576 0.612 ; 
      RECT 3.096 0.252 3.168 0.324 ; 
      RECT 2.88 0.54 2.952 0.612 ; 
      RECT 2.664 0.54 2.736 0.612 ; 
      RECT 2.448 0.252 2.52 0.324 ; 
      RECT 2.232 0.396 2.304 0.468 ; 
      RECT 1.944 0.252 2.016 0.324 ; 
      RECT 1.784 0.396 1.856 0.468 ; 
      RECT 1.564 0.54 1.636 0.612 ; 
      RECT 1.26 0.252 1.332 0.324 ; 
      RECT 0.804 0.252 0.876 0.324 ; 
      RECT 0.612 0.54 0.684 0.612 ; 
      RECT 0.064 0.54 0.136 0.612 ; 
  END 
END DFFLQNx1_ASAP7_6t_SL 


MACRO DFFLQNx2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFFLQNx2_ASAP7_6t_SL 0 0 ; 
  SIZE 4.536 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.704 0.756 ; 
        RECT 0.376 0.108 0.704 0.18 ; 
        RECT 0.288 0.28 0.468 0.352 ; 
        RECT 0.376 0.108 0.468 0.352 ; 
        RECT 0.376 0.532 0.46 0.756 ; 
        RECT 0.288 0.532 0.46 0.604 ; 
        RECT 0.288 0.28 0.36 0.604 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.08 0.684 1.568 0.756 ; 
        RECT 1.004 0.108 1.352 0.18 ; 
        RECT 1.08 0.108 1.152 0.756 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 3.812 0.684 4.248 0.756 ; 
        RECT 4.176 0.108 4.248 0.756 ; 
        RECT 3.812 0.108 4.248 0.18 ; 
    END 
  END QN 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 4.536 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.536 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 3.448 0.54 3.596 0.612 ; 
      RECT 3.524 0.36 3.596 0.612 ; 
      RECT 3.236 0.684 3.512 0.756 ; 
      RECT 3.236 0.512 3.312 0.756 ; 
      RECT 3.24 0.108 3.312 0.756 ; 
      RECT 3.076 0.512 3.312 0.584 ; 
      RECT 3.24 0.108 3.512 0.18 ; 
      RECT 2.536 0.684 2.952 0.756 ; 
      RECT 2.88 0.112 2.952 0.756 ; 
      RECT 2.752 0.112 2.952 0.184 ; 
      RECT 2.616 0.54 2.776 0.612 ; 
      RECT 2.664 0.372 2.736 0.612 ; 
      RECT 2.448 0.252 2.52 0.488 ; 
      RECT 2.404 0.252 2.56 0.324 ; 
      RECT 2.088 0.604 2.412 0.676 ; 
      RECT 2.088 0.108 2.16 0.676 ; 
      RECT 1.976 0.484 2.16 0.556 ; 
      RECT 2.088 0.108 2.512 0.18 ; 
      RECT 1.692 0.684 1.856 0.756 ; 
      RECT 1.784 0.108 1.856 0.756 ; 
      RECT 1.476 0.108 1.856 0.18 ; 
      RECT 1.508 0.54 1.656 0.612 ; 
      RECT 1.584 0.36 1.656 0.612 ; 
      RECT 1.224 0.396 1.472 0.468 ; 
      RECT 1.224 0.252 1.296 0.468 ; 
      RECT 1.224 0.252 1.508 0.324 ; 
      RECT 0.828 0.684 0.976 0.756 ; 
      RECT 0.9 0.344 0.976 0.756 ; 
      RECT 0.804 0.344 0.976 0.416 ; 
      RECT 0.804 0.232 0.876 0.416 ; 
      RECT 0.572 0.54 0.732 0.612 ; 
      RECT 0.572 0.396 0.644 0.612 ; 
      RECT 0.064 0.684 0.252 0.756 ; 
      RECT 0.064 0.108 0.136 0.756 ; 
      RECT 0.064 0.108 0.272 0.18 ; 
      RECT 3.096 0.176 3.168 0.412 ; 
      RECT 2.232 0.288 2.304 0.488 ; 
      RECT 1.944 0.176 2.016 0.36 ; 
    LAYER M2 ; 
      RECT 2.88 0.54 3.596 0.612 ; 
      RECT 0.784 0.252 3.188 0.324 ; 
      RECT 0.064 0.54 2.736 0.612 ; 
      RECT 1.784 0.396 2.304 0.468 ; 
    LAYER V1 ; 
      RECT 3.504 0.54 3.576 0.612 ; 
      RECT 3.096 0.252 3.168 0.324 ; 
      RECT 2.88 0.54 2.952 0.612 ; 
      RECT 2.664 0.54 2.736 0.612 ; 
      RECT 2.448 0.252 2.52 0.324 ; 
      RECT 2.232 0.396 2.304 0.468 ; 
      RECT 1.944 0.252 2.016 0.324 ; 
      RECT 1.784 0.396 1.856 0.468 ; 
      RECT 1.564 0.54 1.636 0.612 ; 
      RECT 1.26 0.252 1.332 0.324 ; 
      RECT 0.804 0.252 0.876 0.324 ; 
      RECT 0.612 0.54 0.684 0.612 ; 
      RECT 0.064 0.54 0.136 0.612 ; 
  END 
END DFFLQNx2_ASAP7_6t_SL 


MACRO DFFLQNx3_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFFLQNx3_ASAP7_6t_SL 0 0 ; 
  SIZE 4.752 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.704 0.756 ; 
        RECT 0.376 0.108 0.704 0.18 ; 
        RECT 0.288 0.28 0.468 0.352 ; 
        RECT 0.376 0.108 0.468 0.352 ; 
        RECT 0.376 0.532 0.46 0.756 ; 
        RECT 0.288 0.532 0.46 0.604 ; 
        RECT 0.288 0.28 0.36 0.604 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.08 0.684 1.568 0.756 ; 
        RECT 1.004 0.108 1.352 0.18 ; 
        RECT 1.08 0.108 1.152 0.756 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.028 0.684 4.676 0.756 ; 
        RECT 4.604 0.108 4.676 0.756 ; 
        RECT 4.044 0.108 4.676 0.18 ; 
    END 
  END QN 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 4.752 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.752 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 3.448 0.54 3.596 0.612 ; 
      RECT 3.524 0.36 3.596 0.612 ; 
      RECT 3.236 0.684 3.512 0.756 ; 
      RECT 3.236 0.512 3.312 0.756 ; 
      RECT 3.24 0.108 3.312 0.756 ; 
      RECT 3.076 0.512 3.312 0.584 ; 
      RECT 3.24 0.108 3.512 0.18 ; 
      RECT 2.536 0.684 2.952 0.756 ; 
      RECT 2.88 0.112 2.952 0.756 ; 
      RECT 2.752 0.112 2.952 0.184 ; 
      RECT 2.616 0.54 2.776 0.612 ; 
      RECT 2.664 0.372 2.736 0.612 ; 
      RECT 2.448 0.252 2.52 0.488 ; 
      RECT 2.404 0.252 2.56 0.324 ; 
      RECT 2.088 0.604 2.412 0.676 ; 
      RECT 2.088 0.108 2.16 0.676 ; 
      RECT 1.976 0.484 2.16 0.556 ; 
      RECT 2.088 0.108 2.512 0.18 ; 
      RECT 1.692 0.684 1.856 0.756 ; 
      RECT 1.784 0.108 1.856 0.756 ; 
      RECT 1.476 0.108 1.856 0.18 ; 
      RECT 1.508 0.54 1.656 0.612 ; 
      RECT 1.584 0.36 1.656 0.612 ; 
      RECT 1.224 0.396 1.472 0.468 ; 
      RECT 1.224 0.252 1.296 0.468 ; 
      RECT 1.224 0.252 1.508 0.324 ; 
      RECT 0.828 0.684 0.976 0.756 ; 
      RECT 0.9 0.344 0.976 0.756 ; 
      RECT 0.804 0.344 0.976 0.416 ; 
      RECT 0.804 0.232 0.876 0.416 ; 
      RECT 0.572 0.54 0.732 0.612 ; 
      RECT 0.572 0.396 0.644 0.612 ; 
      RECT 0.064 0.684 0.252 0.756 ; 
      RECT 0.064 0.108 0.136 0.756 ; 
      RECT 0.064 0.108 0.272 0.18 ; 
      RECT 3.096 0.176 3.168 0.412 ; 
      RECT 2.232 0.288 2.304 0.488 ; 
      RECT 1.944 0.176 2.016 0.36 ; 
    LAYER M2 ; 
      RECT 2.88 0.54 3.596 0.612 ; 
      RECT 0.784 0.252 3.188 0.324 ; 
      RECT 0.064 0.54 2.736 0.612 ; 
      RECT 1.784 0.396 2.304 0.468 ; 
    LAYER V1 ; 
      RECT 3.504 0.54 3.576 0.612 ; 
      RECT 3.096 0.252 3.168 0.324 ; 
      RECT 2.88 0.54 2.952 0.612 ; 
      RECT 2.664 0.54 2.736 0.612 ; 
      RECT 2.448 0.252 2.52 0.324 ; 
      RECT 2.232 0.396 2.304 0.468 ; 
      RECT 1.944 0.252 2.016 0.324 ; 
      RECT 1.784 0.396 1.856 0.468 ; 
      RECT 1.564 0.54 1.636 0.612 ; 
      RECT 1.26 0.252 1.332 0.324 ; 
      RECT 0.804 0.252 0.876 0.324 ; 
      RECT 0.612 0.54 0.684 0.612 ; 
      RECT 0.064 0.54 0.136 0.612 ; 
  END 
END DFFLQNx3_ASAP7_6t_SL 


MACRO DFFLQx4_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFFLQx4_ASAP7_6t_SL 0 0 ; 
  SIZE 5.4 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.704 0.756 ; 
        RECT 0.376 0.108 0.704 0.18 ; 
        RECT 0.288 0.28 0.468 0.352 ; 
        RECT 0.376 0.108 0.468 0.352 ; 
        RECT 0.376 0.532 0.46 0.756 ; 
        RECT 0.288 0.532 0.46 0.604 ; 
        RECT 0.288 0.28 0.36 0.604 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.08 0.684 1.568 0.756 ; 
        RECT 1.004 0.108 1.352 0.18 ; 
        RECT 1.08 0.108 1.152 0.756 ; 
    END 
  END D 
  PIN Q 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.5 0.684 5.332 0.756 ; 
        RECT 5.252 0.108 5.332 0.756 ; 
        RECT 4.5 0.108 5.332 0.18 ; 
        RECT 4.5 0.588 4.572 0.756 ; 
        RECT 4.5 0.108 4.572 0.276 ; 
    END 
  END Q 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 5.4 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.4 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 4.048 0.684 4.392 0.756 ; 
      RECT 4.32 0.108 4.392 0.756 ; 
      RECT 4.32 0.392 4.7 0.464 ; 
      RECT 4.048 0.108 4.392 0.18 ; 
      RECT 3.448 0.54 3.596 0.612 ; 
      RECT 3.524 0.36 3.596 0.612 ; 
      RECT 3.236 0.684 3.512 0.756 ; 
      RECT 3.236 0.512 3.312 0.756 ; 
      RECT 3.24 0.108 3.312 0.756 ; 
      RECT 3.076 0.512 3.312 0.584 ; 
      RECT 3.24 0.108 3.512 0.18 ; 
      RECT 2.536 0.684 2.952 0.756 ; 
      RECT 2.88 0.112 2.952 0.756 ; 
      RECT 2.752 0.112 2.952 0.184 ; 
      RECT 2.616 0.54 2.776 0.612 ; 
      RECT 2.664 0.372 2.736 0.612 ; 
      RECT 2.448 0.252 2.52 0.488 ; 
      RECT 2.404 0.252 2.56 0.324 ; 
      RECT 2.088 0.604 2.412 0.676 ; 
      RECT 2.088 0.108 2.16 0.676 ; 
      RECT 1.976 0.484 2.16 0.556 ; 
      RECT 2.088 0.108 2.512 0.18 ; 
      RECT 1.692 0.684 1.856 0.756 ; 
      RECT 1.784 0.108 1.856 0.756 ; 
      RECT 1.476 0.108 1.856 0.18 ; 
      RECT 1.508 0.54 1.656 0.612 ; 
      RECT 1.584 0.36 1.656 0.612 ; 
      RECT 1.224 0.396 1.472 0.468 ; 
      RECT 1.224 0.252 1.296 0.468 ; 
      RECT 1.224 0.252 1.508 0.324 ; 
      RECT 0.828 0.684 0.976 0.756 ; 
      RECT 0.9 0.344 0.976 0.756 ; 
      RECT 0.804 0.344 0.976 0.416 ; 
      RECT 0.804 0.232 0.876 0.416 ; 
      RECT 0.572 0.54 0.732 0.612 ; 
      RECT 0.572 0.396 0.644 0.612 ; 
      RECT 0.064 0.684 0.252 0.756 ; 
      RECT 0.064 0.108 0.136 0.756 ; 
      RECT 0.064 0.108 0.272 0.18 ; 
      RECT 3.096 0.176 3.168 0.412 ; 
      RECT 2.232 0.288 2.304 0.488 ; 
      RECT 1.944 0.176 2.016 0.36 ; 
    LAYER M2 ; 
      RECT 2.88 0.54 3.596 0.612 ; 
      RECT 0.784 0.252 3.188 0.324 ; 
      RECT 0.064 0.54 2.736 0.612 ; 
      RECT 1.784 0.396 2.304 0.468 ; 
    LAYER V1 ; 
      RECT 3.504 0.54 3.576 0.612 ; 
      RECT 3.096 0.252 3.168 0.324 ; 
      RECT 2.88 0.54 2.952 0.612 ; 
      RECT 2.664 0.54 2.736 0.612 ; 
      RECT 2.448 0.252 2.52 0.324 ; 
      RECT 2.232 0.396 2.304 0.468 ; 
      RECT 1.944 0.252 2.016 0.324 ; 
      RECT 1.784 0.396 1.856 0.468 ; 
      RECT 1.564 0.54 1.636 0.612 ; 
      RECT 1.26 0.252 1.332 0.324 ; 
      RECT 0.804 0.252 0.876 0.324 ; 
      RECT 0.612 0.54 0.684 0.612 ; 
      RECT 0.064 0.54 0.136 0.612 ; 
  END 
END DFFLQx4_ASAP7_6t_SL 


MACRO DHLx1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DHLx1_ASAP7_6t_SL 0 0 ; 
  SIZE 3.24 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.704 0.756 ; 
        RECT 0.376 0.108 0.704 0.18 ; 
        RECT 0.288 0.26 0.468 0.332 ; 
        RECT 0.376 0.108 0.468 0.332 ; 
        RECT 0.376 0.512 0.448 0.756 ; 
        RECT 0.288 0.512 0.448 0.584 ; 
        RECT 0.288 0.26 0.36 0.584 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.08 0.684 1.352 0.756 ; 
        RECT 1.08 0.108 1.352 0.18 ; 
        RECT 1.08 0.396 1.224 0.468 ; 
        RECT 1.08 0.108 1.152 0.756 ; 
    END 
  END D 
  PIN Q 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.744 0.684 3.168 0.756 ; 
        RECT 3.096 0.108 3.168 0.756 ; 
        RECT 2.744 0.108 3.168 0.18 ; 
    END 
  END Q 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.24 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.24 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.32 0.684 2.628 0.756 ; 
      RECT 2.556 0.108 2.628 0.756 ; 
      RECT 2.016 0.28 2.208 0.352 ; 
      RECT 2.136 0.108 2.208 0.352 ; 
      RECT 2.136 0.108 2.628 0.18 ; 
      RECT 2.412 0.252 2.484 0.504 ; 
      RECT 2.308 0.252 2.484 0.324 ; 
      RECT 1.476 0.684 1.872 0.756 ; 
      RECT 1.8 0.108 1.872 0.756 ; 
      RECT 1.652 0.108 1.872 0.18 ; 
      RECT 1.584 0.252 1.656 0.504 ; 
      RECT 1.528 0.252 1.696 0.324 ; 
      RECT 1.352 0.54 1.5 0.612 ; 
      RECT 1.368 0.34 1.44 0.612 ; 
      RECT 0.828 0.684 0.98 0.756 ; 
      RECT 0.908 0.108 0.98 0.756 ; 
      RECT 0.828 0.108 0.98 0.18 ; 
      RECT 0.572 0.54 0.792 0.612 ; 
      RECT 0.72 0.396 0.792 0.612 ; 
      RECT 0.552 0.396 0.792 0.468 ; 
      RECT 0.064 0.684 0.272 0.756 ; 
      RECT 0.064 0.108 0.136 0.756 ; 
      RECT 0.064 0.108 0.272 0.18 ; 
      RECT 2.016 0.452 2.088 0.688 ; 
    LAYER M2 ; 
      RECT 1.8 0.252 2.44 0.324 ; 
      RECT 0.064 0.54 2.108 0.612 ; 
      RECT 0.888 0.252 1.656 0.324 ; 
    LAYER V1 ; 
      RECT 2.34 0.252 2.412 0.324 ; 
      RECT 2.016 0.54 2.088 0.612 ; 
      RECT 1.8 0.252 1.872 0.324 ; 
      RECT 1.584 0.252 1.656 0.324 ; 
      RECT 1.368 0.54 1.44 0.612 ; 
      RECT 0.908 0.252 0.98 0.324 ; 
      RECT 0.612 0.54 0.684 0.612 ; 
      RECT 0.064 0.54 0.136 0.612 ; 
  END 
END DHLx1_ASAP7_6t_SL 


MACRO DHLx2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DHLx2_ASAP7_6t_SL 0 0 ; 
  SIZE 3.456 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.704 0.756 ; 
        RECT 0.376 0.108 0.704 0.18 ; 
        RECT 0.288 0.26 0.468 0.332 ; 
        RECT 0.376 0.108 0.468 0.332 ; 
        RECT 0.376 0.512 0.448 0.756 ; 
        RECT 0.288 0.512 0.448 0.584 ; 
        RECT 0.288 0.26 0.36 0.584 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.08 0.684 1.352 0.756 ; 
        RECT 1.08 0.108 1.352 0.18 ; 
        RECT 1.08 0.396 1.224 0.468 ; 
        RECT 1.08 0.108 1.152 0.756 ; 
    END 
  END D 
  PIN Q 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.752 0.684 3.168 0.756 ; 
        RECT 3.096 0.108 3.168 0.756 ; 
        RECT 2.752 0.108 3.168 0.18 ; 
    END 
  END Q 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.456 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.456 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.32 0.684 2.628 0.756 ; 
      RECT 2.556 0.108 2.628 0.756 ; 
      RECT 2.016 0.28 2.208 0.352 ; 
      RECT 2.136 0.108 2.208 0.352 ; 
      RECT 2.136 0.108 2.628 0.18 ; 
      RECT 2.412 0.252 2.484 0.504 ; 
      RECT 2.308 0.252 2.484 0.324 ; 
      RECT 1.476 0.684 1.872 0.756 ; 
      RECT 1.8 0.108 1.872 0.756 ; 
      RECT 1.652 0.108 1.872 0.18 ; 
      RECT 1.584 0.252 1.656 0.504 ; 
      RECT 1.528 0.252 1.696 0.324 ; 
      RECT 1.352 0.54 1.5 0.612 ; 
      RECT 1.368 0.34 1.44 0.612 ; 
      RECT 0.828 0.684 0.98 0.756 ; 
      RECT 0.908 0.108 0.98 0.756 ; 
      RECT 0.828 0.108 0.98 0.18 ; 
      RECT 0.572 0.54 0.792 0.612 ; 
      RECT 0.72 0.396 0.792 0.612 ; 
      RECT 0.552 0.396 0.792 0.468 ; 
      RECT 0.064 0.684 0.272 0.756 ; 
      RECT 0.064 0.108 0.136 0.756 ; 
      RECT 0.064 0.108 0.272 0.18 ; 
      RECT 2.016 0.452 2.088 0.688 ; 
    LAYER M2 ; 
      RECT 1.8 0.252 2.44 0.324 ; 
      RECT 0.064 0.54 2.108 0.612 ; 
      RECT 0.888 0.252 1.656 0.324 ; 
    LAYER V1 ; 
      RECT 2.34 0.252 2.412 0.324 ; 
      RECT 2.016 0.54 2.088 0.612 ; 
      RECT 1.8 0.252 1.872 0.324 ; 
      RECT 1.584 0.252 1.656 0.324 ; 
      RECT 1.368 0.54 1.44 0.612 ; 
      RECT 0.908 0.252 0.98 0.324 ; 
      RECT 0.612 0.54 0.684 0.612 ; 
      RECT 0.064 0.54 0.136 0.612 ; 
  END 
END DHLx2_ASAP7_6t_SL 


MACRO DHLx3_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DHLx3_ASAP7_6t_SL 0 0 ; 
  SIZE 3.672 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.704 0.756 ; 
        RECT 0.376 0.108 0.704 0.18 ; 
        RECT 0.288 0.26 0.468 0.332 ; 
        RECT 0.376 0.108 0.468 0.332 ; 
        RECT 0.376 0.512 0.448 0.756 ; 
        RECT 0.288 0.512 0.448 0.584 ; 
        RECT 0.288 0.26 0.36 0.584 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.08 0.684 1.352 0.756 ; 
        RECT 1.08 0.108 1.352 0.18 ; 
        RECT 1.08 0.396 1.224 0.468 ; 
        RECT 1.08 0.108 1.152 0.756 ; 
    END 
  END D 
  PIN Q 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.896 0.684 3.524 0.756 ; 
        RECT 2.908 0.108 3.524 0.18 ; 
        RECT 3.096 0.108 3.168 0.756 ; 
    END 
  END Q 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.672 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.672 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.32 0.684 2.628 0.756 ; 
      RECT 2.556 0.108 2.628 0.756 ; 
      RECT 2.016 0.28 2.208 0.352 ; 
      RECT 2.136 0.108 2.208 0.352 ; 
      RECT 2.136 0.108 2.628 0.18 ; 
      RECT 2.412 0.252 2.484 0.504 ; 
      RECT 2.308 0.252 2.484 0.324 ; 
      RECT 1.476 0.684 1.872 0.756 ; 
      RECT 1.8 0.108 1.872 0.756 ; 
      RECT 1.652 0.108 1.872 0.18 ; 
      RECT 1.584 0.252 1.656 0.504 ; 
      RECT 1.528 0.252 1.696 0.324 ; 
      RECT 1.352 0.54 1.5 0.612 ; 
      RECT 1.368 0.34 1.44 0.612 ; 
      RECT 0.828 0.684 0.98 0.756 ; 
      RECT 0.908 0.108 0.98 0.756 ; 
      RECT 0.828 0.108 0.98 0.18 ; 
      RECT 0.572 0.54 0.792 0.612 ; 
      RECT 0.72 0.396 0.792 0.612 ; 
      RECT 0.552 0.396 0.792 0.468 ; 
      RECT 0.064 0.684 0.272 0.756 ; 
      RECT 0.064 0.108 0.136 0.756 ; 
      RECT 0.064 0.108 0.272 0.18 ; 
      RECT 2.016 0.452 2.088 0.688 ; 
    LAYER M2 ; 
      RECT 1.8 0.252 2.44 0.324 ; 
      RECT 0.064 0.54 2.108 0.612 ; 
      RECT 0.888 0.252 1.656 0.324 ; 
    LAYER V1 ; 
      RECT 2.34 0.252 2.412 0.324 ; 
      RECT 2.016 0.54 2.088 0.612 ; 
      RECT 1.8 0.252 1.872 0.324 ; 
      RECT 1.584 0.252 1.656 0.324 ; 
      RECT 1.368 0.54 1.44 0.612 ; 
      RECT 0.908 0.252 0.98 0.324 ; 
      RECT 0.612 0.54 0.684 0.612 ; 
      RECT 0.064 0.54 0.136 0.612 ; 
  END 
END DHLx3_ASAP7_6t_SL 


MACRO DLLx1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DLLx1_ASAP7_6t_SL 0 0 ; 
  SIZE 3.24 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.704 0.756 ; 
        RECT 0.376 0.108 0.704 0.18 ; 
        RECT 0.376 0.532 0.468 0.756 ; 
        RECT 0.288 0.28 0.448 0.352 ; 
        RECT 0.376 0.108 0.448 0.352 ; 
        RECT 0.288 0.532 0.468 0.604 ; 
        RECT 0.288 0.28 0.36 0.604 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.08 0.684 1.352 0.756 ; 
        RECT 1.08 0.108 1.352 0.18 ; 
        RECT 1.08 0.396 1.224 0.468 ; 
        RECT 1.08 0.108 1.152 0.756 ; 
    END 
  END D 
  PIN Q 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.744 0.684 3.168 0.756 ; 
        RECT 3.096 0.108 3.168 0.756 ; 
        RECT 2.744 0.108 3.168 0.18 ; 
    END 
  END Q 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.24 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.24 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.136 0.684 2.628 0.756 ; 
      RECT 2.556 0.108 2.628 0.756 ; 
      RECT 2.136 0.512 2.208 0.756 ; 
      RECT 2.016 0.512 2.208 0.584 ; 
      RECT 2.32 0.108 2.628 0.18 ; 
      RECT 2.308 0.54 2.484 0.612 ; 
      RECT 2.412 0.36 2.484 0.612 ; 
      RECT 1.652 0.684 1.872 0.756 ; 
      RECT 1.8 0.108 1.872 0.756 ; 
      RECT 1.476 0.108 1.872 0.18 ; 
      RECT 1.528 0.54 1.696 0.612 ; 
      RECT 1.584 0.36 1.656 0.612 ; 
      RECT 1.368 0.252 1.44 0.524 ; 
      RECT 1.352 0.252 1.5 0.324 ; 
      RECT 0.828 0.684 0.98 0.756 ; 
      RECT 0.908 0.108 0.98 0.756 ; 
      RECT 0.828 0.108 0.98 0.18 ; 
      RECT 0.552 0.396 0.792 0.468 ; 
      RECT 0.72 0.252 0.792 0.468 ; 
      RECT 0.572 0.252 0.792 0.324 ; 
      RECT 0.064 0.684 0.272 0.756 ; 
      RECT 0.064 0.108 0.136 0.756 ; 
      RECT 0.064 0.108 0.272 0.18 ; 
      RECT 2.016 0.176 2.088 0.412 ; 
    LAYER M2 ; 
      RECT 1.8 0.54 2.44 0.612 ; 
      RECT 0.064 0.252 2.108 0.324 ; 
      RECT 0.888 0.54 1.656 0.612 ; 
    LAYER V1 ; 
      RECT 2.34 0.54 2.412 0.612 ; 
      RECT 2.016 0.252 2.088 0.324 ; 
      RECT 1.8 0.54 1.872 0.612 ; 
      RECT 1.584 0.54 1.656 0.612 ; 
      RECT 1.368 0.252 1.44 0.324 ; 
      RECT 0.908 0.54 0.98 0.612 ; 
      RECT 0.612 0.252 0.684 0.324 ; 
      RECT 0.064 0.252 0.136 0.324 ; 
  END 
END DLLx1_ASAP7_6t_SL 


MACRO DLLx2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DLLx2_ASAP7_6t_SL 0 0 ; 
  SIZE 3.456 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.704 0.756 ; 
        RECT 0.376 0.108 0.704 0.18 ; 
        RECT 0.376 0.532 0.468 0.756 ; 
        RECT 0.288 0.28 0.448 0.352 ; 
        RECT 0.376 0.108 0.448 0.352 ; 
        RECT 0.288 0.532 0.468 0.604 ; 
        RECT 0.288 0.28 0.36 0.604 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.08 0.684 1.352 0.756 ; 
        RECT 1.08 0.108 1.352 0.18 ; 
        RECT 1.08 0.396 1.224 0.468 ; 
        RECT 1.08 0.108 1.152 0.756 ; 
    END 
  END D 
  PIN Q 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.744 0.684 3.168 0.756 ; 
        RECT 3.096 0.108 3.168 0.756 ; 
        RECT 2.744 0.108 3.168 0.18 ; 
    END 
  END Q 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.456 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.456 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.136 0.684 2.628 0.756 ; 
      RECT 2.556 0.108 2.628 0.756 ; 
      RECT 2.136 0.512 2.208 0.756 ; 
      RECT 2.016 0.512 2.208 0.584 ; 
      RECT 2.32 0.108 2.628 0.18 ; 
      RECT 2.308 0.54 2.484 0.612 ; 
      RECT 2.412 0.36 2.484 0.612 ; 
      RECT 1.652 0.684 1.872 0.756 ; 
      RECT 1.8 0.108 1.872 0.756 ; 
      RECT 1.476 0.108 1.872 0.18 ; 
      RECT 1.528 0.54 1.696 0.612 ; 
      RECT 1.584 0.36 1.656 0.612 ; 
      RECT 1.368 0.252 1.44 0.524 ; 
      RECT 1.352 0.252 1.5 0.324 ; 
      RECT 0.828 0.684 0.98 0.756 ; 
      RECT 0.908 0.108 0.98 0.756 ; 
      RECT 0.828 0.108 0.98 0.18 ; 
      RECT 0.552 0.396 0.792 0.468 ; 
      RECT 0.72 0.252 0.792 0.468 ; 
      RECT 0.572 0.252 0.792 0.324 ; 
      RECT 0.064 0.684 0.272 0.756 ; 
      RECT 0.064 0.108 0.136 0.756 ; 
      RECT 0.064 0.108 0.272 0.18 ; 
      RECT 2.016 0.176 2.088 0.412 ; 
    LAYER M2 ; 
      RECT 1.8 0.54 2.44 0.612 ; 
      RECT 0.064 0.252 2.108 0.324 ; 
      RECT 0.888 0.54 1.656 0.612 ; 
    LAYER V1 ; 
      RECT 2.34 0.54 2.412 0.612 ; 
      RECT 2.016 0.252 2.088 0.324 ; 
      RECT 1.8 0.54 1.872 0.612 ; 
      RECT 1.584 0.54 1.656 0.612 ; 
      RECT 1.368 0.252 1.44 0.324 ; 
      RECT 0.908 0.54 0.98 0.612 ; 
      RECT 0.612 0.252 0.684 0.324 ; 
      RECT 0.064 0.252 0.136 0.324 ; 
  END 
END DLLx2_ASAP7_6t_SL 


MACRO DLLx3_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DLLx3_ASAP7_6t_SL 0 0 ; 
  SIZE 3.672 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.704 0.756 ; 
        RECT 0.376 0.108 0.704 0.18 ; 
        RECT 0.376 0.532 0.468 0.756 ; 
        RECT 0.288 0.28 0.448 0.352 ; 
        RECT 0.376 0.108 0.448 0.352 ; 
        RECT 0.288 0.532 0.468 0.604 ; 
        RECT 0.288 0.28 0.36 0.604 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.08 0.684 1.352 0.756 ; 
        RECT 1.08 0.108 1.352 0.18 ; 
        RECT 1.08 0.396 1.224 0.468 ; 
        RECT 1.08 0.108 1.152 0.756 ; 
    END 
  END D 
  PIN Q 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.908 0.684 3.524 0.756 ; 
        RECT 2.892 0.108 3.524 0.18 ; 
        RECT 3.096 0.108 3.168 0.756 ; 
    END 
  END Q 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.672 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.672 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.136 0.684 2.628 0.756 ; 
      RECT 2.556 0.108 2.628 0.756 ; 
      RECT 2.136 0.512 2.208 0.756 ; 
      RECT 2.016 0.512 2.208 0.584 ; 
      RECT 2.32 0.108 2.628 0.18 ; 
      RECT 2.308 0.54 2.484 0.612 ; 
      RECT 2.412 0.36 2.484 0.612 ; 
      RECT 1.652 0.684 1.872 0.756 ; 
      RECT 1.8 0.108 1.872 0.756 ; 
      RECT 1.476 0.108 1.872 0.18 ; 
      RECT 1.528 0.54 1.696 0.612 ; 
      RECT 1.584 0.36 1.656 0.612 ; 
      RECT 1.368 0.252 1.44 0.524 ; 
      RECT 1.352 0.252 1.5 0.324 ; 
      RECT 0.828 0.684 0.98 0.756 ; 
      RECT 0.908 0.108 0.98 0.756 ; 
      RECT 0.828 0.108 0.98 0.18 ; 
      RECT 0.552 0.396 0.792 0.468 ; 
      RECT 0.72 0.252 0.792 0.468 ; 
      RECT 0.572 0.252 0.792 0.324 ; 
      RECT 0.064 0.684 0.272 0.756 ; 
      RECT 0.064 0.108 0.136 0.756 ; 
      RECT 0.064 0.108 0.272 0.18 ; 
      RECT 2.016 0.176 2.088 0.412 ; 
    LAYER M2 ; 
      RECT 1.8 0.54 2.44 0.612 ; 
      RECT 0.064 0.252 2.108 0.324 ; 
      RECT 0.888 0.54 1.656 0.612 ; 
    LAYER V1 ; 
      RECT 2.34 0.54 2.412 0.612 ; 
      RECT 2.016 0.252 2.088 0.324 ; 
      RECT 1.8 0.54 1.872 0.612 ; 
      RECT 1.584 0.54 1.656 0.612 ; 
      RECT 1.368 0.252 1.44 0.324 ; 
      RECT 0.908 0.54 0.98 0.612 ; 
      RECT 0.612 0.252 0.684 0.324 ; 
      RECT 0.064 0.252 0.136 0.324 ; 
  END 
END DLLx3_ASAP7_6t_SL 


MACRO FAxp33_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FAxp33_ASAP7_6t_SL 0 0 ; 
  SIZE 3.024 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.024 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.024 0.036 ; 
    END 
  END VSS 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.448 0.252 2.596 0.324 ; 
        RECT 2.448 0.252 2.52 0.5 ; 
        RECT 1.556 0.396 1.724 0.468 ; 
        RECT 1.652 0.232 1.724 0.468 ; 
        RECT 0.072 0.252 0.312 0.324 ; 
        RECT 0.072 0.252 0.144 0.52 ; 
      LAYER M2 ; 
        RECT 0.16 0.252 2.572 0.324 ; 
      LAYER V1 ; 
        RECT 0.18 0.252 0.252 0.324 ; 
        RECT 1.652 0.252 1.724 0.324 ; 
        RECT 2.472 0.252 2.544 0.324 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.744 0.684 2.952 0.756 ; 
        RECT 2.88 0.352 2.952 0.756 ; 
        RECT 1.24 0.684 1.46 0.756 ; 
        RECT 1.24 0.376 1.312 0.756 ; 
        RECT 0.72 0.54 1.312 0.612 ; 
        RECT 0.72 0.376 0.792 0.612 ; 
      LAYER M2 ; 
        RECT 1.24 0.684 2.868 0.756 ; 
      LAYER V1 ; 
        RECT 1.26 0.684 1.332 0.756 ; 
        RECT 2.772 0.684 2.844 0.756 ; 
    END 
  END B 
  PIN CI 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.172 0.396 2.344 0.468 ; 
        RECT 2.172 0.316 2.244 0.5 ; 
        RECT 1.8 0.368 1.872 0.58 ; 
        RECT 0.948 0.396 1.168 0.468 ; 
        RECT 1.096 0.252 1.168 0.468 ; 
        RECT 0.948 0.252 1.168 0.324 ; 
      LAYER M2 ; 
        RECT 0.9 0.396 2.36 0.468 ; 
      LAYER V1 ; 
        RECT 1.008 0.396 1.08 0.468 ; 
        RECT 1.8 0.396 1.872 0.468 ; 
        RECT 2.256 0.396 2.328 0.468 ; 
    END 
  END CI 
  PIN CON 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.004 0.288 2.076 0.54 ; 
        RECT 1.944 0.468 2.016 0.688 ; 
        RECT 0.496 0.152 0.832 0.224 ; 
        RECT 0.56 0.54 0.632 0.704 ; 
        RECT 0.496 0.152 0.568 0.612 ; 
      LAYER M2 ; 
        RECT 0.504 0.54 2.036 0.612 ; 
      LAYER V1 ; 
        RECT 0.536 0.54 0.608 0.612 ; 
        RECT 1.944 0.54 2.016 0.612 ; 
    END 
  END CON 
  PIN SN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.384 0.54 1.672 0.612 ; 
        RECT 1.384 0.108 1.568 0.18 ; 
        RECT 1.384 0.108 1.456 0.612 ; 
      LAYER M2 ; 
        RECT 1.452 0.108 2.596 0.18 ; 
      LAYER V1 ; 
        RECT 1.476 0.108 1.548 0.18 ; 
    END 
  END SN 
  OBS 
    LAYER M1 ; 
      RECT 2.124 0.108 2.648 0.18 ; 
      RECT 2.156 0.612 2.596 0.684 ; 
      RECT 0.972 0.108 1.18 0.18 ; 
      RECT 0.78 0.684 1.116 0.756 ; 
      RECT 0.16 0.684 0.348 0.756 ; 
      RECT 0.16 0.108 0.328 0.18 ; 
    LAYER M2 ; 
      RECT 0.16 0.108 1.136 0.18 ; 
      RECT 0.16 0.684 0.924 0.756 ; 
    LAYER V1 ; 
      RECT 1.044 0.108 1.116 0.18 ; 
      RECT 0.828 0.684 0.9 0.756 ; 
      RECT 0.18 0.108 0.252 0.18 ; 
      RECT 0.18 0.684 0.252 0.756 ; 
  END 
END FAxp33_ASAP7_6t_SL 


MACRO FILLER_ASAP7_6t_SL 
  CLASS CORE SPACER ; 
  ORIGIN 0 0 ; 
  FOREIGN FILLER_ASAP7_6t_SL 0 0 ; 
  SIZE 0.432 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 0.432 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.432 0.036 ; 
    END 
  END VSS 
END FILLER_ASAP7_6t_SL 


MACRO FILLERxp5_ASAP7_6t_SL 
  CLASS CORE SPACER ; 
  ORIGIN 0 0 ; 
  FOREIGN FILLERxp5_ASAP7_6t_SL 0 0 ; 
  SIZE 0.216 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 0.216 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.216 0.036 ; 
    END 
  END VSS 
END FILLERxp5_ASAP7_6t_SL 


MACRO HAxp5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN HAxp5_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.676 0.396 1.44 0.468 ; 
        RECT 0.676 0.108 0.748 0.468 ; 
        RECT 0.072 0.108 0.748 0.18 ; 
        RECT 0.072 0.684 0.272 0.756 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.28 0.396 0.576 0.468 ; 
        RECT 0.28 0.252 0.576 0.324 ; 
        RECT 0.352 0.54 0.572 0.612 ; 
        RECT 0.352 0.396 0.424 0.612 ; 
        RECT 0.28 0.252 0.352 0.468 ; 
    END 
  END B 
  PIN CON 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.704 0.54 1.656 0.612 ; 
        RECT 1.584 0.252 1.656 0.612 ; 
        RECT 0.848 0.252 1.656 0.324 ; 
        RECT 0.396 0.684 0.776 0.756 ; 
        RECT 0.704 0.54 0.776 0.756 ; 
    END 
  END CON 
  PIN SN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.684 1.88 0.756 ; 
        RECT 1.808 0.108 1.88 0.756 ; 
        RECT 1.692 0.108 1.88 0.18 ; 
    END 
  END SN 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 1.044 0.108 1.548 0.18 ; 
  END 
END HAxp5_ASAP7_6t_SL 


MACRO HB1x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN HB1x1_ASAP7_6t_SL 0 0 ; 
  SIZE 0.864 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.54 0.292 0.612 ; 
        RECT 0.072 0.396 0.292 0.468 ; 
        RECT 0.072 0.252 0.292 0.324 ; 
        RECT 0.072 0.252 0.144 0.612 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 0.864 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.864 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.684 0.792 0.756 ; 
        RECT 0.72 0.108 0.792 0.756 ; 
        RECT 0.592 0.108 0.792 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.144 0.684 0.476 0.756 ; 
      RECT 0.404 0.108 0.476 0.756 ; 
      RECT 0.404 0.396 0.596 0.468 ; 
      RECT 0.136 0.108 0.476 0.18 ; 
  END 
END HB1x1_ASAP7_6t_SL 


MACRO HB2x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN HB2x1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.08 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.38 0.468 ; 
        RECT 0.072 0.684 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.08 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.08 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.684 1.008 0.756 ; 
        RECT 0.936 0.108 1.008 0.756 ; 
        RECT 0.808 0.108 1.008 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.396 0.684 0.576 0.756 ; 
      RECT 0.504 0.108 0.576 0.756 ; 
      RECT 0.504 0.396 0.812 0.468 ; 
      RECT 0.396 0.108 0.576 0.18 ; 
  END 
END HB2x1_ASAP7_6t_SL 


MACRO HB3x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN HB3x1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.38 0.468 ; 
        RECT 0.072 0.684 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.684 1.224 0.756 ; 
        RECT 1.152 0.108 1.224 0.756 ; 
        RECT 1.024 0.108 1.224 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.396 0.684 0.792 0.756 ; 
      RECT 0.72 0.108 0.792 0.756 ; 
      RECT 0.72 0.396 1.028 0.468 ; 
      RECT 0.396 0.108 0.792 0.18 ; 
  END 
END HB3x1_ASAP7_6t_SL 


MACRO HB4x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN HB4x1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.064 0.396 0.404 0.468 ; 
        RECT 0.064 0.684 0.272 0.756 ; 
        RECT 0.064 0.108 0.272 0.18 ; 
        RECT 0.064 0.108 0.136 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.24 0.684 1.44 0.756 ; 
        RECT 1.368 0.108 1.44 0.756 ; 
        RECT 1.24 0.108 1.44 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.396 0.684 0.792 0.756 ; 
      RECT 0.72 0.108 0.792 0.756 ; 
      RECT 0.72 0.396 1.244 0.468 ; 
      RECT 0.396 0.108 0.792 0.18 ; 
  END 
END HB4x1_ASAP7_6t_SL 


MACRO ICGx10_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ICGx10_ASAP7_6t_SL 0 0 ; 
  SIZE 6.696 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 3.72 0.54 3.944 0.612 ; 
        RECT 3.872 0.44 3.944 0.612 ; 
        RECT 2.448 0.54 3.04 0.612 ; 
        RECT 2.968 0.44 3.04 0.612 ; 
        RECT 2.596 0.108 2.824 0.18 ; 
        RECT 2.448 0.252 2.668 0.324 ; 
        RECT 2.596 0.108 2.668 0.324 ; 
        RECT 2.448 0.252 2.52 0.612 ; 
        RECT 1.584 0.452 1.656 0.688 ; 
        RECT 0.92 0.54 1.068 0.612 ; 
        RECT 0.936 0.34 1.008 0.612 ; 
      LAYER M2 ; 
        RECT 0.9 0.54 3.832 0.612 ; 
      LAYER V1 ; 
        RECT 0.936 0.54 1.008 0.612 ; 
        RECT 1.584 0.54 1.656 0.612 ; 
        RECT 2.672 0.54 2.744 0.612 ; 
        RECT 3.76 0.54 3.832 0.612 ; 
    END 
  END CLK 
  PIN ENA 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.392 0.36 0.464 ; 
        RECT 0.072 0.684 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END ENA 
  PIN GCLK 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.392 0.684 6.524 0.756 ; 
        RECT 6.444 0.108 6.524 0.756 ; 
        RECT 4.404 0.108 6.524 0.18 ; 
    END 
  END GCLK 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.54 0.576 0.612 ; 
        RECT 0.504 0.252 0.576 0.612 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END SE 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 6.696 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 6.696 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.74 0.684 4.248 0.756 ; 
      RECT 4.176 0.54 4.248 0.756 ; 
      RECT 4.176 0.54 4.464 0.612 ; 
      RECT 4.392 0.252 4.464 0.612 ; 
      RECT 4.192 0.252 4.464 0.324 ; 
      RECT 4.192 0.108 4.264 0.324 ; 
      RECT 2.988 0.108 4.264 0.18 ; 
      RECT 3.148 0.396 3.408 0.468 ; 
      RECT 2.628 0.396 2.86 0.468 ; 
      RECT 2.788 0.252 2.86 0.468 ; 
      RECT 3.148 0.252 3.22 0.468 ; 
      RECT 2.788 0.252 3.22 0.324 ; 
      RECT 2.236 0.684 2.556 0.756 ; 
      RECT 2.236 0.108 2.308 0.756 ; 
      RECT 2.236 0.108 2.412 0.18 ; 
      RECT 1.888 0.684 2.136 0.756 ; 
      RECT 2.064 0.108 2.136 0.756 ; 
      RECT 1.584 0.28 1.776 0.352 ; 
      RECT 1.704 0.108 1.776 0.352 ; 
      RECT 1.704 0.108 2.136 0.18 ; 
      RECT 1.024 0.684 1.44 0.756 ; 
      RECT 1.368 0.108 1.44 0.756 ; 
      RECT 1.22 0.108 1.44 0.18 ; 
      RECT 1.152 0.252 1.224 0.504 ; 
      RECT 1.096 0.252 1.264 0.324 ; 
      RECT 0.396 0.684 0.792 0.756 ; 
      RECT 0.72 0.108 0.792 0.756 ; 
      RECT 0.396 0.108 0.792 0.18 ; 
      RECT 4.076 0.396 4.292 0.468 ; 
      RECT 1.848 0.28 1.92 0.504 ; 
    LAYER M2 ; 
      RECT 1.32 0.396 4.28 0.468 ; 
      RECT 1.128 0.252 2.344 0.324 ; 
    LAYER V1 ; 
      RECT 4.168 0.396 4.24 0.468 ; 
      RECT 2.672 0.396 2.744 0.468 ; 
      RECT 2.236 0.252 2.308 0.324 ; 
      RECT 1.848 0.396 1.92 0.468 ; 
      RECT 1.368 0.396 1.44 0.468 ; 
      RECT 1.152 0.252 1.224 0.324 ; 
  END 
END ICGx10_ASAP7_6t_SL 


MACRO ICGx12_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ICGx12_ASAP7_6t_SL 0 0 ; 
  SIZE 7.128 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 3.72 0.54 3.944 0.612 ; 
        RECT 3.872 0.44 3.944 0.612 ; 
        RECT 2.448 0.54 3.04 0.612 ; 
        RECT 2.968 0.44 3.04 0.612 ; 
        RECT 2.596 0.108 2.824 0.18 ; 
        RECT 2.448 0.252 2.668 0.324 ; 
        RECT 2.596 0.108 2.668 0.324 ; 
        RECT 2.448 0.252 2.52 0.612 ; 
        RECT 1.584 0.452 1.656 0.688 ; 
        RECT 0.92 0.54 1.068 0.612 ; 
        RECT 0.936 0.34 1.008 0.612 ; 
      LAYER M2 ; 
        RECT 0.9 0.54 3.832 0.612 ; 
      LAYER V1 ; 
        RECT 0.936 0.54 1.008 0.612 ; 
        RECT 1.584 0.54 1.656 0.612 ; 
        RECT 2.672 0.54 2.744 0.612 ; 
        RECT 3.76 0.54 3.832 0.612 ; 
    END 
  END CLK 
  PIN ENA 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.216 0.392 0.36 0.464 ; 
        RECT 0.14 0.54 0.288 0.612 ; 
        RECT 0.216 0.108 0.288 0.612 ; 
        RECT 0.14 0.108 0.288 0.18 ; 
    END 
  END ENA 
  PIN GCLK 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.38 0.684 6.884 0.756 ; 
        RECT 6.812 0.108 6.884 0.756 ; 
        RECT 4.392 0.108 6.884 0.18 ; 
    END 
  END GCLK 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.54 0.576 0.612 ; 
        RECT 0.504 0.252 0.576 0.612 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END SE 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 7.128 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 7.128 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.74 0.684 4.248 0.756 ; 
      RECT 4.176 0.54 4.248 0.756 ; 
      RECT 4.176 0.54 4.464 0.612 ; 
      RECT 4.392 0.252 4.464 0.612 ; 
      RECT 4.192 0.252 4.464 0.324 ; 
      RECT 4.192 0.108 4.264 0.324 ; 
      RECT 2.988 0.108 4.264 0.18 ; 
      RECT 3.148 0.396 3.408 0.468 ; 
      RECT 2.628 0.396 2.86 0.468 ; 
      RECT 2.788 0.252 2.86 0.468 ; 
      RECT 3.148 0.252 3.22 0.468 ; 
      RECT 2.788 0.252 3.22 0.324 ; 
      RECT 2.236 0.684 2.556 0.756 ; 
      RECT 2.236 0.108 2.308 0.756 ; 
      RECT 2.236 0.108 2.412 0.18 ; 
      RECT 1.888 0.684 2.136 0.756 ; 
      RECT 2.064 0.108 2.136 0.756 ; 
      RECT 1.584 0.28 1.776 0.352 ; 
      RECT 1.704 0.108 1.776 0.352 ; 
      RECT 1.704 0.108 2.136 0.18 ; 
      RECT 1.024 0.684 1.44 0.756 ; 
      RECT 1.368 0.108 1.44 0.756 ; 
      RECT 1.22 0.108 1.44 0.18 ; 
      RECT 1.152 0.252 1.224 0.504 ; 
      RECT 1.096 0.252 1.264 0.324 ; 
      RECT 0.148 0.684 0.792 0.756 ; 
      RECT 0.72 0.108 0.792 0.756 ; 
      RECT 0.396 0.108 0.792 0.18 ; 
      RECT 4.076 0.396 4.292 0.468 ; 
      RECT 1.848 0.28 1.92 0.504 ; 
    LAYER M2 ; 
      RECT 1.32 0.396 4.28 0.468 ; 
      RECT 1.128 0.252 2.344 0.324 ; 
    LAYER V1 ; 
      RECT 4.168 0.396 4.24 0.468 ; 
      RECT 2.672 0.396 2.744 0.468 ; 
      RECT 2.236 0.252 2.308 0.324 ; 
      RECT 1.848 0.396 1.92 0.468 ; 
      RECT 1.368 0.396 1.44 0.468 ; 
      RECT 1.152 0.252 1.224 0.324 ; 
  END 
END ICGx12_ASAP7_6t_SL 


MACRO ICGx1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ICGx1_ASAP7_6t_SL 0 0 ; 
  SIZE 3.888 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 2.448 0.54 3.04 0.612 ; 
        RECT 2.968 0.44 3.04 0.612 ; 
        RECT 2.596 0.108 2.824 0.18 ; 
        RECT 2.448 0.252 2.668 0.324 ; 
        RECT 2.596 0.108 2.668 0.324 ; 
        RECT 2.448 0.252 2.52 0.612 ; 
        RECT 1.584 0.684 1.784 0.756 ; 
        RECT 1.584 0.452 1.656 0.756 ; 
        RECT 0.936 0.108 1.156 0.18 ; 
        RECT 0.92 0.54 1.068 0.612 ; 
        RECT 0.936 0.108 1.008 0.612 ; 
      LAYER M2 ; 
        RECT 0.9 0.54 2.768 0.612 ; 
      LAYER V1 ; 
        RECT 0.936 0.54 1.008 0.612 ; 
        RECT 1.584 0.54 1.656 0.612 ; 
        RECT 2.672 0.54 2.744 0.612 ; 
    END 
  END CLK 
  PIN ENA 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.216 0.392 0.36 0.464 ; 
        RECT 0.14 0.68 0.288 0.756 ; 
        RECT 0.216 0.108 0.288 0.756 ; 
        RECT 0.14 0.108 0.288 0.18 ; 
    END 
  END ENA 
  PIN GCLK 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 3.512 0.684 3.812 0.756 ; 
        RECT 3.74 0.108 3.812 0.756 ; 
        RECT 3.524 0.108 3.812 0.18 ; 
    END 
  END GCLK 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.54 0.576 0.612 ; 
        RECT 0.504 0.252 0.576 0.612 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END SE 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.888 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.888 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.752 0.684 3.384 0.756 ; 
      RECT 3.312 0.54 3.384 0.756 ; 
      RECT 3.312 0.54 3.6 0.612 ; 
      RECT 3.528 0.252 3.6 0.612 ; 
      RECT 3.328 0.252 3.6 0.324 ; 
      RECT 3.328 0.108 3.4 0.324 ; 
      RECT 2.948 0.108 3.4 0.18 ; 
      RECT 3.148 0.396 3.408 0.468 ; 
      RECT 2.628 0.396 2.86 0.468 ; 
      RECT 2.788 0.252 2.86 0.468 ; 
      RECT 3.148 0.252 3.22 0.468 ; 
      RECT 2.788 0.252 3.22 0.324 ; 
      RECT 2.236 0.684 2.556 0.756 ; 
      RECT 2.236 0.108 2.308 0.756 ; 
      RECT 2.236 0.108 2.412 0.18 ; 
      RECT 1.908 0.684 2.136 0.756 ; 
      RECT 2.064 0.108 2.136 0.756 ; 
      RECT 1.584 0.28 1.776 0.352 ; 
      RECT 1.704 0.108 1.776 0.352 ; 
      RECT 1.704 0.108 2.136 0.18 ; 
      RECT 1.024 0.684 1.44 0.756 ; 
      RECT 1.368 0.136 1.44 0.756 ; 
      RECT 1.152 0.252 1.224 0.504 ; 
      RECT 1.108 0.252 1.264 0.324 ; 
      RECT 0.396 0.684 0.792 0.756 ; 
      RECT 0.72 0.108 0.792 0.756 ; 
      RECT 0.396 0.108 0.792 0.18 ; 
      RECT 1.848 0.28 1.92 0.504 ; 
    LAYER M2 ; 
      RECT 1.32 0.396 2.768 0.468 ; 
      RECT 1.128 0.252 2.344 0.324 ; 
    LAYER V1 ; 
      RECT 2.672 0.396 2.744 0.468 ; 
      RECT 2.236 0.252 2.308 0.324 ; 
      RECT 1.848 0.396 1.92 0.468 ; 
      RECT 1.368 0.396 1.44 0.468 ; 
      RECT 1.152 0.252 1.224 0.324 ; 
  END 
END ICGx1_ASAP7_6t_SL 


MACRO ICGx2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ICGx2_ASAP7_6t_SL 0 0 ; 
  SIZE 4.104 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 2.448 0.54 3.04 0.612 ; 
        RECT 2.968 0.44 3.04 0.612 ; 
        RECT 2.596 0.108 2.824 0.18 ; 
        RECT 2.448 0.252 2.668 0.324 ; 
        RECT 2.596 0.108 2.668 0.324 ; 
        RECT 2.448 0.252 2.52 0.612 ; 
        RECT 1.584 0.68 1.784 0.752 ; 
        RECT 1.584 0.452 1.656 0.752 ; 
        RECT 0.936 0.108 1.156 0.18 ; 
        RECT 0.92 0.54 1.068 0.612 ; 
        RECT 0.936 0.108 1.008 0.612 ; 
      LAYER M2 ; 
        RECT 0.9 0.54 2.768 0.612 ; 
      LAYER V1 ; 
        RECT 0.936 0.54 1.008 0.612 ; 
        RECT 1.584 0.54 1.656 0.612 ; 
        RECT 2.672 0.54 2.744 0.612 ; 
    END 
  END CLK 
  PIN ENA 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.216 0.392 0.36 0.464 ; 
        RECT 0.14 0.684 0.288 0.756 ; 
        RECT 0.216 0.108 0.288 0.756 ; 
        RECT 0.14 0.108 0.288 0.18 ; 
    END 
  END ENA 
  PIN GCLK 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 3.516 0.684 3.816 0.756 ; 
        RECT 3.744 0.108 3.816 0.756 ; 
        RECT 3.528 0.108 3.816 0.18 ; 
    END 
  END GCLK 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.54 0.576 0.612 ; 
        RECT 0.504 0.252 0.576 0.612 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END SE 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 4.104 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.104 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.752 0.684 3.384 0.756 ; 
      RECT 3.312 0.54 3.384 0.756 ; 
      RECT 3.312 0.54 3.6 0.612 ; 
      RECT 3.528 0.252 3.6 0.612 ; 
      RECT 3.328 0.252 3.6 0.324 ; 
      RECT 3.328 0.108 3.4 0.324 ; 
      RECT 2.948 0.108 3.4 0.18 ; 
      RECT 3.148 0.396 3.408 0.468 ; 
      RECT 2.628 0.396 2.86 0.468 ; 
      RECT 2.788 0.252 2.86 0.468 ; 
      RECT 3.148 0.252 3.22 0.468 ; 
      RECT 2.788 0.252 3.22 0.324 ; 
      RECT 2.236 0.684 2.556 0.756 ; 
      RECT 2.236 0.108 2.308 0.756 ; 
      RECT 2.236 0.108 2.412 0.18 ; 
      RECT 1.908 0.684 2.136 0.756 ; 
      RECT 2.064 0.108 2.136 0.756 ; 
      RECT 1.584 0.28 1.776 0.352 ; 
      RECT 1.704 0.108 1.776 0.352 ; 
      RECT 1.704 0.108 2.136 0.18 ; 
      RECT 1.024 0.684 1.44 0.756 ; 
      RECT 1.368 0.136 1.44 0.756 ; 
      RECT 1.152 0.252 1.224 0.504 ; 
      RECT 1.108 0.252 1.264 0.324 ; 
      RECT 0.396 0.684 0.792 0.756 ; 
      RECT 0.72 0.108 0.792 0.756 ; 
      RECT 0.396 0.108 0.792 0.18 ; 
      RECT 1.848 0.28 1.92 0.504 ; 
    LAYER M2 ; 
      RECT 1.32 0.396 2.768 0.468 ; 
      RECT 1.128 0.252 2.344 0.324 ; 
    LAYER V1 ; 
      RECT 2.672 0.396 2.744 0.468 ; 
      RECT 2.236 0.252 2.308 0.324 ; 
      RECT 1.848 0.396 1.92 0.468 ; 
      RECT 1.368 0.396 1.44 0.468 ; 
      RECT 1.152 0.252 1.224 0.324 ; 
  END 
END ICGx2_ASAP7_6t_SL 


MACRO ICGx3_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ICGx3_ASAP7_6t_SL 0 0 ; 
  SIZE 4.32 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 2.448 0.54 3.04 0.612 ; 
        RECT 2.968 0.44 3.04 0.612 ; 
        RECT 2.596 0.108 2.824 0.18 ; 
        RECT 2.448 0.252 2.668 0.324 ; 
        RECT 2.596 0.108 2.668 0.324 ; 
        RECT 2.448 0.252 2.52 0.612 ; 
        RECT 1.584 0.684 1.784 0.756 ; 
        RECT 1.584 0.452 1.656 0.756 ; 
        RECT 0.936 0.108 1.156 0.18 ; 
        RECT 0.92 0.54 1.068 0.612 ; 
        RECT 0.936 0.108 1.008 0.612 ; 
      LAYER M2 ; 
        RECT 0.9 0.54 2.768 0.612 ; 
      LAYER V1 ; 
        RECT 0.936 0.54 1.008 0.612 ; 
        RECT 1.584 0.54 1.656 0.612 ; 
        RECT 2.672 0.54 2.744 0.612 ; 
    END 
  END CLK 
  PIN ENA 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.216 0.392 0.36 0.464 ; 
        RECT 0.14 0.684 0.288 0.756 ; 
        RECT 0.216 0.108 0.288 0.756 ; 
        RECT 0.14 0.108 0.288 0.18 ; 
    END 
  END ENA 
  PIN GCLK 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 3.516 0.684 4.164 0.756 ; 
        RECT 3.528 0.108 4.164 0.18 ; 
        RECT 3.744 0.108 3.816 0.756 ; 
    END 
  END GCLK 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.54 0.576 0.612 ; 
        RECT 0.504 0.252 0.576 0.612 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END SE 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 4.32 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.32 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.752 0.684 3.384 0.756 ; 
      RECT 3.312 0.54 3.384 0.756 ; 
      RECT 3.312 0.54 3.6 0.612 ; 
      RECT 3.528 0.252 3.6 0.612 ; 
      RECT 3.328 0.252 3.6 0.324 ; 
      RECT 3.328 0.108 3.4 0.324 ; 
      RECT 2.948 0.108 3.4 0.18 ; 
      RECT 3.148 0.396 3.408 0.468 ; 
      RECT 2.628 0.396 2.86 0.468 ; 
      RECT 2.788 0.252 2.86 0.468 ; 
      RECT 3.148 0.252 3.22 0.468 ; 
      RECT 2.788 0.252 3.22 0.324 ; 
      RECT 2.236 0.684 2.556 0.756 ; 
      RECT 2.236 0.108 2.308 0.756 ; 
      RECT 2.236 0.108 2.412 0.18 ; 
      RECT 1.908 0.684 2.136 0.756 ; 
      RECT 2.064 0.108 2.136 0.756 ; 
      RECT 1.584 0.28 1.776 0.352 ; 
      RECT 1.704 0.108 1.776 0.352 ; 
      RECT 1.704 0.108 2.136 0.18 ; 
      RECT 1.024 0.684 1.44 0.756 ; 
      RECT 1.368 0.136 1.44 0.756 ; 
      RECT 1.152 0.252 1.224 0.504 ; 
      RECT 1.108 0.252 1.264 0.324 ; 
      RECT 0.396 0.684 0.792 0.756 ; 
      RECT 0.72 0.108 0.792 0.756 ; 
      RECT 0.396 0.108 0.792 0.18 ; 
      RECT 1.848 0.28 1.92 0.504 ; 
    LAYER M2 ; 
      RECT 1.32 0.396 2.768 0.468 ; 
      RECT 1.128 0.252 2.344 0.324 ; 
    LAYER V1 ; 
      RECT 2.672 0.396 2.744 0.468 ; 
      RECT 2.236 0.252 2.308 0.324 ; 
      RECT 1.848 0.396 1.92 0.468 ; 
      RECT 1.368 0.396 1.44 0.468 ; 
      RECT 1.152 0.252 1.224 0.324 ; 
  END 
END ICGx3_ASAP7_6t_SL 


MACRO ICGx4_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ICGx4_ASAP7_6t_SL 0 0 ; 
  SIZE 5.4 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 3.72 0.54 3.944 0.612 ; 
        RECT 3.872 0.44 3.944 0.612 ; 
        RECT 2.448 0.54 3.04 0.612 ; 
        RECT 2.968 0.44 3.04 0.612 ; 
        RECT 2.596 0.108 2.824 0.18 ; 
        RECT 2.448 0.252 2.668 0.324 ; 
        RECT 2.596 0.108 2.668 0.324 ; 
        RECT 2.448 0.252 2.52 0.612 ; 
        RECT 1.584 0.684 1.784 0.756 ; 
        RECT 1.584 0.452 1.656 0.756 ; 
        RECT 0.932 0.108 1.168 0.18 ; 
        RECT 0.92 0.54 1.068 0.612 ; 
        RECT 0.936 0.108 1.008 0.612 ; 
      LAYER M2 ; 
        RECT 0.9 0.54 3.832 0.612 ; 
      LAYER V1 ; 
        RECT 0.936 0.54 1.008 0.612 ; 
        RECT 1.584 0.54 1.656 0.612 ; 
        RECT 2.672 0.54 2.744 0.612 ; 
        RECT 3.76 0.54 3.832 0.612 ; 
    END 
  END CLK 
  PIN ENA 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.216 0.392 0.36 0.464 ; 
        RECT 0.14 0.684 0.288 0.756 ; 
        RECT 0.216 0.108 0.288 0.756 ; 
        RECT 0.14 0.108 0.288 0.18 ; 
    END 
  END ENA 
  PIN GCLK 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.38 0.684 5.176 0.756 ; 
        RECT 5.104 0.108 5.176 0.756 ; 
        RECT 4.392 0.108 5.176 0.18 ; 
    END 
  END GCLK 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.54 0.576 0.612 ; 
        RECT 0.504 0.252 0.576 0.612 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END SE 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 5.4 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.4 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.74 0.684 4.248 0.756 ; 
      RECT 4.176 0.54 4.248 0.756 ; 
      RECT 4.176 0.54 4.464 0.612 ; 
      RECT 4.392 0.252 4.464 0.612 ; 
      RECT 4.192 0.252 4.464 0.324 ; 
      RECT 4.192 0.108 4.264 0.324 ; 
      RECT 2.988 0.108 4.264 0.18 ; 
      RECT 3.148 0.396 3.408 0.468 ; 
      RECT 2.628 0.396 2.86 0.468 ; 
      RECT 2.788 0.252 2.86 0.468 ; 
      RECT 3.148 0.252 3.22 0.468 ; 
      RECT 2.788 0.252 3.22 0.324 ; 
      RECT 2.236 0.684 2.556 0.756 ; 
      RECT 2.236 0.108 2.308 0.756 ; 
      RECT 2.236 0.108 2.412 0.18 ; 
      RECT 1.908 0.684 2.136 0.756 ; 
      RECT 2.064 0.108 2.136 0.756 ; 
      RECT 1.584 0.28 1.776 0.352 ; 
      RECT 1.704 0.108 1.776 0.352 ; 
      RECT 1.704 0.108 2.136 0.18 ; 
      RECT 1.024 0.684 1.44 0.756 ; 
      RECT 1.368 0.136 1.44 0.756 ; 
      RECT 1.152 0.252 1.224 0.504 ; 
      RECT 1.108 0.252 1.264 0.324 ; 
      RECT 0.396 0.684 0.792 0.756 ; 
      RECT 0.72 0.108 0.792 0.756 ; 
      RECT 0.396 0.108 0.792 0.18 ; 
      RECT 4.076 0.396 4.292 0.468 ; 
      RECT 1.848 0.28 1.92 0.504 ; 
    LAYER M2 ; 
      RECT 1.32 0.396 4.28 0.468 ; 
      RECT 1.128 0.252 2.344 0.324 ; 
    LAYER V1 ; 
      RECT 4.168 0.396 4.24 0.468 ; 
      RECT 2.672 0.396 2.744 0.468 ; 
      RECT 2.236 0.252 2.308 0.324 ; 
      RECT 1.848 0.396 1.92 0.468 ; 
      RECT 1.368 0.396 1.44 0.468 ; 
      RECT 1.152 0.252 1.224 0.324 ; 
  END 
END ICGx4_ASAP7_6t_SL 


MACRO ICGx5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ICGx5_ASAP7_6t_SL 0 0 ; 
  SIZE 5.616 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 3.72 0.54 3.944 0.612 ; 
        RECT 3.872 0.44 3.944 0.612 ; 
        RECT 2.448 0.54 3.04 0.612 ; 
        RECT 2.968 0.44 3.04 0.612 ; 
        RECT 2.596 0.108 2.824 0.18 ; 
        RECT 2.448 0.252 2.668 0.324 ; 
        RECT 2.596 0.108 2.668 0.324 ; 
        RECT 2.448 0.252 2.52 0.612 ; 
        RECT 1.584 0.684 1.784 0.756 ; 
        RECT 1.584 0.452 1.656 0.756 ; 
        RECT 0.936 0.108 1.156 0.18 ; 
        RECT 0.92 0.54 1.068 0.612 ; 
        RECT 0.936 0.108 1.008 0.612 ; 
      LAYER M2 ; 
        RECT 0.9 0.54 3.832 0.612 ; 
      LAYER V1 ; 
        RECT 0.936 0.54 1.008 0.612 ; 
        RECT 1.584 0.54 1.656 0.612 ; 
        RECT 2.672 0.54 2.744 0.612 ; 
        RECT 3.76 0.54 3.832 0.612 ; 
    END 
  END CLK 
  PIN ENA 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.216 0.392 0.36 0.464 ; 
        RECT 0.14 0.68 0.288 0.756 ; 
        RECT 0.216 0.108 0.288 0.756 ; 
        RECT 0.14 0.108 0.288 0.18 ; 
    END 
  END ENA 
  PIN GCLK 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.38 0.684 5.528 0.756 ; 
        RECT 5.456 0.108 5.528 0.756 ; 
        RECT 4.392 0.108 5.528 0.18 ; 
    END 
  END GCLK 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.54 0.576 0.612 ; 
        RECT 0.504 0.252 0.576 0.612 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END SE 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 5.616 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.616 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.74 0.684 4.248 0.756 ; 
      RECT 4.176 0.54 4.248 0.756 ; 
      RECT 4.176 0.54 4.464 0.612 ; 
      RECT 4.392 0.252 4.464 0.612 ; 
      RECT 4.192 0.252 4.464 0.324 ; 
      RECT 4.192 0.108 4.264 0.324 ; 
      RECT 2.988 0.108 4.264 0.18 ; 
      RECT 3.148 0.396 3.408 0.468 ; 
      RECT 2.628 0.396 2.86 0.468 ; 
      RECT 2.788 0.252 2.86 0.468 ; 
      RECT 3.148 0.252 3.22 0.468 ; 
      RECT 2.788 0.252 3.22 0.324 ; 
      RECT 2.236 0.684 2.556 0.756 ; 
      RECT 2.236 0.108 2.308 0.756 ; 
      RECT 2.236 0.108 2.412 0.18 ; 
      RECT 1.908 0.684 2.136 0.756 ; 
      RECT 2.064 0.108 2.136 0.756 ; 
      RECT 1.584 0.28 1.776 0.352 ; 
      RECT 1.704 0.108 1.776 0.352 ; 
      RECT 1.704 0.108 2.136 0.18 ; 
      RECT 1.024 0.684 1.44 0.756 ; 
      RECT 1.368 0.136 1.44 0.756 ; 
      RECT 1.152 0.252 1.224 0.504 ; 
      RECT 1.108 0.252 1.264 0.324 ; 
      RECT 0.396 0.684 0.792 0.756 ; 
      RECT 0.72 0.108 0.792 0.756 ; 
      RECT 0.396 0.108 0.792 0.18 ; 
      RECT 4.076 0.396 4.292 0.468 ; 
      RECT 1.848 0.28 1.92 0.504 ; 
    LAYER M2 ; 
      RECT 1.32 0.396 4.28 0.468 ; 
      RECT 1.128 0.252 2.344 0.324 ; 
    LAYER V1 ; 
      RECT 4.168 0.396 4.24 0.468 ; 
      RECT 2.672 0.396 2.744 0.468 ; 
      RECT 2.236 0.252 2.308 0.324 ; 
      RECT 1.848 0.396 1.92 0.468 ; 
      RECT 1.368 0.396 1.44 0.468 ; 
      RECT 1.152 0.252 1.224 0.324 ; 
  END 
END ICGx5_ASAP7_6t_SL 


MACRO ICGx8_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ICGx8_ASAP7_6t_SL 0 0 ; 
  SIZE 6.264 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 3.72 0.54 3.944 0.612 ; 
        RECT 3.872 0.44 3.944 0.612 ; 
        RECT 2.448 0.54 3.04 0.612 ; 
        RECT 2.968 0.44 3.04 0.612 ; 
        RECT 2.596 0.108 2.864 0.18 ; 
        RECT 2.448 0.252 2.668 0.324 ; 
        RECT 2.596 0.108 2.668 0.324 ; 
        RECT 2.448 0.252 2.52 0.612 ; 
        RECT 1.584 0.452 1.656 0.688 ; 
        RECT 0.92 0.54 1.068 0.612 ; 
        RECT 0.936 0.34 1.008 0.612 ; 
      LAYER M2 ; 
        RECT 0.9 0.54 3.832 0.612 ; 
      LAYER V1 ; 
        RECT 0.936 0.54 1.008 0.612 ; 
        RECT 1.584 0.54 1.656 0.612 ; 
        RECT 2.672 0.54 2.744 0.612 ; 
        RECT 3.76 0.54 3.832 0.612 ; 
    END 
  END CLK 
  PIN ENA 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.392 0.38 0.464 ; 
        RECT 0.072 0.684 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END ENA 
  PIN GCLK 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.48 0.684 6.032 0.756 ; 
        RECT 5.96 0.108 6.032 0.756 ; 
        RECT 4.48 0.108 6.032 0.18 ; 
    END 
  END GCLK 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.54 0.576 0.612 ; 
        RECT 0.504 0.252 0.576 0.612 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END SE 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 6.264 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 6.264 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.74 0.684 4.248 0.756 ; 
      RECT 4.176 0.54 4.248 0.756 ; 
      RECT 4.176 0.54 4.436 0.612 ; 
      RECT 4.364 0.252 4.436 0.612 ; 
      RECT 4.364 0.4 5.456 0.472 ; 
      RECT 4.192 0.252 4.436 0.324 ; 
      RECT 4.192 0.108 4.264 0.324 ; 
      RECT 2.988 0.108 4.264 0.18 ; 
      RECT 3.148 0.396 3.408 0.468 ; 
      RECT 2.628 0.396 2.86 0.468 ; 
      RECT 2.788 0.252 2.86 0.468 ; 
      RECT 3.148 0.252 3.22 0.468 ; 
      RECT 2.788 0.252 3.22 0.324 ; 
      RECT 2.208 0.684 2.412 0.756 ; 
      RECT 2.208 0.108 2.28 0.756 ; 
      RECT 2.208 0.108 2.412 0.18 ; 
      RECT 1.888 0.684 2.136 0.756 ; 
      RECT 2.064 0.108 2.136 0.756 ; 
      RECT 1.584 0.28 1.776 0.352 ; 
      RECT 1.704 0.108 1.776 0.352 ; 
      RECT 1.704 0.108 2.136 0.18 ; 
      RECT 1.024 0.684 1.44 0.756 ; 
      RECT 1.368 0.108 1.44 0.756 ; 
      RECT 1.22 0.108 1.44 0.18 ; 
      RECT 1.152 0.252 1.224 0.504 ; 
      RECT 1.096 0.252 1.264 0.324 ; 
      RECT 0.396 0.684 0.792 0.756 ; 
      RECT 0.72 0.108 0.792 0.756 ; 
      RECT 0.396 0.108 0.792 0.18 ; 
      RECT 4.076 0.396 4.264 0.468 ; 
      RECT 1.848 0.28 1.92 0.504 ; 
    LAYER M2 ; 
      RECT 1.32 0.396 4.28 0.468 ; 
      RECT 1.132 0.252 2.3 0.324 ; 
    LAYER V1 ; 
      RECT 4.168 0.396 4.24 0.468 ; 
      RECT 2.672 0.396 2.744 0.468 ; 
      RECT 2.208 0.252 2.28 0.324 ; 
      RECT 1.848 0.396 1.92 0.468 ; 
      RECT 1.368 0.396 1.44 0.468 ; 
      RECT 1.152 0.252 1.224 0.324 ; 
  END 
END ICGx8_ASAP7_6t_SL 


MACRO INVx11_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx11_ASAP7_6t_SL 0 0 ; 
  SIZE 2.808 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.312 0.468 ; 
        RECT 0.072 0.608 0.276 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.808 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.808 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 2.736 0.756 ; 
        RECT 2.664 0.108 2.736 0.756 ; 
        RECT 0.376 0.108 2.736 0.18 ; 
    END 
  END Y 
END INVx11_ASAP7_6t_SL 


MACRO INVx13_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx13_ASAP7_6t_SL 0 0 ; 
  SIZE 3.24 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.312 0.468 ; 
        RECT 0.072 0.684 0.22 0.756 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.24 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.24 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 3.168 0.756 ; 
        RECT 3.096 0.108 3.168 0.756 ; 
        RECT 0.376 0.108 3.168 0.18 ; 
    END 
  END Y 
END INVx13_ASAP7_6t_SL 


MACRO INVx1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx1_ASAP7_6t_SL 0 0 ; 
  SIZE 0.648 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.312 0.468 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 0.648 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.648 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.576 0.756 ; 
        RECT 0.504 0.108 0.576 0.756 ; 
        RECT 0.376 0.108 0.576 0.18 ; 
    END 
  END Y 
END INVx1_ASAP7_6t_SL 


MACRO INVx2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx2_ASAP7_6t_SL 0 0 ; 
  SIZE 0.864 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 0.864 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.864 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.792 0.756 ; 
        RECT 0.72 0.108 0.792 0.756 ; 
        RECT 0.376 0.108 0.792 0.18 ; 
    END 
  END Y 
END INVx2_ASAP7_6t_SL 


MACRO INVx3_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx3_ASAP7_6t_SL 0 0 ; 
  SIZE 1.08 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.312 0.468 ; 
        RECT 0.072 0.608 0.276 0.756 ; 
        RECT 0.072 0.108 0.276 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.08 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.08 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 1.008 0.756 ; 
        RECT 0.936 0.108 1.008 0.756 ; 
        RECT 0.376 0.108 1.008 0.18 ; 
    END 
  END Y 
END INVx3_ASAP7_6t_SL 


MACRO INVx4_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx4_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.312 0.468 ; 
        RECT 0.072 0.684 0.22 0.756 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 1.224 0.756 ; 
        RECT 1.152 0.108 1.224 0.756 ; 
        RECT 0.376 0.108 1.224 0.18 ; 
    END 
  END Y 
END INVx4_ASAP7_6t_SL 


MACRO INVx5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx5_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.38 0.468 ; 
        RECT 0.072 0.684 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.684 1.44 0.756 ; 
        RECT 1.368 0.108 1.44 0.756 ; 
        RECT 0.396 0.108 1.44 0.18 ; 
    END 
  END Y 
END INVx5_ASAP7_6t_SL 


MACRO INVx6_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx6_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.312 0.468 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 1.656 0.756 ; 
        RECT 1.584 0.108 1.656 0.756 ; 
        RECT 0.376 0.108 1.656 0.18 ; 
    END 
  END Y 
END INVx6_ASAP7_6t_SL 


MACRO INVx8_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx8_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.312 0.468 ; 
        RECT 0.072 0.608 0.276 0.756 ; 
        RECT 0.072 0.108 0.276 0.288 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 2.088 0.756 ; 
        RECT 2.016 0.108 2.088 0.756 ; 
        RECT 0.376 0.108 2.088 0.18 ; 
    END 
  END Y 
END INVx8_ASAP7_6t_SL 


MACRO INVxp5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVxp5_ASAP7_6t_SL 0 0 ; 
  SIZE 0.648 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.312 0.468 ; 
        RECT 0.072 0.684 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 0.648 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.648 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.684 0.576 0.756 ; 
        RECT 0.504 0.108 0.576 0.756 ; 
        RECT 0.396 0.108 0.576 0.18 ; 
    END 
  END Y 
END INVxp5_ASAP7_6t_SL 


MACRO MAJIxp5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MAJIxp5_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.216 0.396 0.712 0.468 ; 
        RECT 0.14 0.684 0.288 0.756 ; 
        RECT 0.216 0.396 0.288 0.756 ; 
    END 
  END A 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.164 0.54 1.608 0.612 ; 
        RECT 1.164 0.252 1.404 0.324 ; 
        RECT 1.164 0.252 1.236 0.612 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.684 1.612 0.756 ; 
        RECT 0.58 0.108 1.332 0.18 ; 
        RECT 1.02 0.108 1.092 0.756 ; 
    END 
  END Y 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.16 0.108 1.572 0.18 ; 
      LAYER M1 ; 
        RECT 1.544 0.396 1.692 0.468 ; 
        RECT 1.62 0.108 1.692 0.468 ; 
        RECT 1.456 0.108 1.692 0.18 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.108 0.144 0.492 ; 
      LAYER V1 ; 
        RECT 0.18 0.108 0.252 0.18 ; 
        RECT 1.476 0.108 1.548 0.18 ; 
    END 
  END B 
  OBS 
    LAYER M1 ; 
      RECT 0.372 0.252 0.92 0.324 ; 
      RECT 0.396 0.54 0.92 0.612 ; 
  END 
END MAJIxp5_ASAP7_6t_SL 


MACRO MAJx1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MAJx1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.508 0.54 0.728 0.612 ; 
        RECT 0.656 0.252 0.728 0.612 ; 
        RECT 0.508 0.252 0.728 0.324 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.684 1.428 0.756 ; 
        RECT 1.356 0.36 1.428 0.756 ; 
        RECT 0.072 0.252 0.224 0.324 ; 
        RECT 0.072 0.252 0.144 0.756 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.828 0.54 1.008 0.612 ; 
        RECT 0.936 0.252 1.008 0.612 ; 
        RECT 0.828 0.252 1.008 0.324 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.672 0.684 1.872 0.756 ; 
        RECT 1.8 0.108 1.872 0.756 ; 
        RECT 1.672 0.108 1.872 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.12 0.54 1.284 0.612 ; 
      RECT 1.212 0.108 1.284 0.612 ; 
      RECT 0.244 0.54 0.408 0.612 ; 
      RECT 0.336 0.108 0.408 0.612 ; 
      RECT 1.5 0.396 1.648 0.468 ; 
      RECT 1.5 0.108 1.572 0.468 ; 
      RECT 0.112 0.108 1.572 0.18 ; 
  END 
END MAJx1_ASAP7_6t_SL 


MACRO MAJx2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MAJx2_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.508 0.54 0.728 0.612 ; 
        RECT 0.656 0.252 0.728 0.612 ; 
        RECT 0.508 0.252 0.728 0.324 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.684 1.428 0.756 ; 
        RECT 1.356 0.36 1.428 0.756 ; 
        RECT 0.072 0.252 0.224 0.324 ; 
        RECT 0.072 0.252 0.144 0.756 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.828 0.54 1.008 0.612 ; 
        RECT 0.936 0.252 1.008 0.612 ; 
        RECT 0.828 0.252 1.008 0.324 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.672 0.684 1.872 0.756 ; 
        RECT 1.8 0.108 1.872 0.756 ; 
        RECT 1.672 0.108 1.872 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.12 0.54 1.284 0.612 ; 
      RECT 1.212 0.108 1.284 0.612 ; 
      RECT 0.244 0.54 0.408 0.612 ; 
      RECT 0.336 0.108 0.408 0.612 ; 
      RECT 1.5 0.396 1.648 0.468 ; 
      RECT 1.5 0.108 1.572 0.468 ; 
      RECT 0.112 0.108 1.572 0.18 ; 
  END 
END MAJx2_ASAP7_6t_SL 


MACRO MAJx3_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MAJx3_ASAP7_6t_SL 0 0 ; 
  SIZE 2.376 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.508 0.54 0.728 0.612 ; 
        RECT 0.656 0.252 0.728 0.612 ; 
        RECT 0.508 0.252 0.728 0.324 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.684 1.428 0.756 ; 
        RECT 1.356 0.36 1.428 0.756 ; 
        RECT 0.072 0.252 0.224 0.324 ; 
        RECT 0.072 0.252 0.144 0.756 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.828 0.54 1.008 0.612 ; 
        RECT 0.936 0.252 1.008 0.612 ; 
        RECT 0.828 0.252 1.008 0.324 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.376 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.672 0.684 2.22 0.756 ; 
        RECT 1.672 0.108 2.22 0.18 ; 
        RECT 1.8 0.108 1.872 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.12 0.54 1.284 0.612 ; 
      RECT 1.212 0.108 1.284 0.612 ; 
      RECT 0.244 0.54 0.408 0.612 ; 
      RECT 0.336 0.108 0.408 0.612 ; 
      RECT 1.5 0.396 1.648 0.468 ; 
      RECT 1.5 0.108 1.572 0.468 ; 
      RECT 0.112 0.108 1.572 0.18 ; 
  END 
END MAJx3_ASAP7_6t_SL 


MACRO NAND2x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND2x1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.336 0.468 ; 
        RECT 0.072 0.252 0.292 0.324 ; 
        RECT 0.072 0.684 0.272 0.756 ; 
        RECT 0.072 0.252 0.144 0.756 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.46 0.396 0.92 0.468 ; 
        RECT 0.46 0.54 0.68 0.612 ; 
        RECT 0.46 0.252 0.68 0.324 ; 
        RECT 0.46 0.252 0.532 0.612 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.684 1.244 0.756 ; 
        RECT 1.172 0.252 1.244 0.756 ; 
        RECT 0.808 0.252 1.244 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.108 1.136 0.18 ; 
  END 
END NAND2x1_ASAP7_6t_SL 


MACRO NAND2x1p5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND2x1p5_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.336 0.468 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.468 0.54 1.352 0.612 ; 
        RECT 0.468 0.396 1.136 0.468 ; 
        RECT 0.468 0.252 0.688 0.324 ; 
        RECT 0.468 0.252 0.54 0.612 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 1.656 0.756 ; 
        RECT 1.584 0.108 1.656 0.756 ; 
        RECT 1.044 0.108 1.656 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.828 0.252 1.352 0.324 ; 
      RECT 0.376 0.108 0.92 0.18 ; 
  END 
END NAND2x1p5_ASAP7_6t_SL 


MACRO NAND2x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND2x2_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.968 0.54 1.188 0.612 ; 
        RECT 1.116 0.396 1.188 0.612 ; 
        RECT 0.968 0.396 1.188 0.468 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.652 0.54 1.872 0.612 ; 
        RECT 1.8 0.396 1.872 0.612 ; 
        RECT 1.288 0.396 1.872 0.468 ; 
        RECT 1.288 0.252 1.36 0.468 ; 
        RECT 0.728 0.252 1.36 0.324 ; 
        RECT 0.288 0.396 0.8 0.468 ; 
        RECT 0.728 0.252 0.8 0.468 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.684 2.088 0.756 ; 
        RECT 2.016 0.252 2.088 0.756 ; 
        RECT 1.672 0.252 2.088 0.324 ; 
        RECT 0.072 0.252 0.488 0.324 ; 
        RECT 0.072 0.252 0.144 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.108 2 0.18 ; 
  END 
END NAND2x2_ASAP7_6t_SL 


MACRO NAND2xp5R_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND2xp5R_ASAP7_6t_SL 0 0 ; 
  SIZE 0.864 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.124 0.684 0.272 0.756 ; 
        RECT 0.2 0.108 0.272 0.756 ; 
        RECT 0.124 0.108 0.272 0.18 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.42 0.54 0.64 0.612 ; 
        RECT 0.42 0.396 0.64 0.468 ; 
        RECT 0.42 0.108 0.492 0.612 ; 
        RECT 0.344 0.108 0.492 0.256 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 0.864 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.864 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.828 0.756 ; 
        RECT 0.756 0.108 0.828 0.756 ; 
        RECT 0.592 0.108 0.828 0.18 ; 
    END 
  END Y 
END NAND2xp5R_ASAP7_6t_SL 


MACRO NAND2xp5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND2xp5_ASAP7_6t_SL 0 0 ; 
  SIZE 0.864 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.068 0.684 0.272 0.756 ; 
        RECT 0.068 0.108 0.272 0.256 ; 
        RECT 0.068 0.108 0.14 0.756 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.356 0.396 0.576 0.468 ; 
        RECT 0.356 0.108 0.504 0.612 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 0.864 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.864 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.684 0.792 0.756 ; 
        RECT 0.72 0.108 0.792 0.756 ; 
        RECT 0.592 0.108 0.792 0.256 ; 
    END 
  END Y 
END NAND2xp5_ASAP7_6t_SL 


MACRO NAND3x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND3x1_ASAP7_6t_SL 0 0 ; 
  SIZE 2.376 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.484 0.54 1.812 0.612 ; 
        RECT 1.484 0.396 1.808 0.468 ; 
        RECT 1.484 0.396 1.556 0.612 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.512 0.396 1.352 0.468 ; 
        RECT 0.512 0.252 0.788 0.324 ; 
        RECT 0.512 0.592 0.708 0.756 ; 
        RECT 0.512 0.252 0.584 0.756 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.336 0.468 ; 
        RECT 0.072 0.684 0.32 0.756 ; 
        RECT 0.072 0.108 0.272 0.28 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.376 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.684 2.304 0.756 ; 
        RECT 2.232 0.108 2.304 0.756 ; 
        RECT 1.672 0.108 2.304 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.024 0.252 2 0.324 ; 
      RECT 0.376 0.108 1.352 0.18 ; 
  END 
END NAND3x1_ASAP7_6t_SL 


MACRO NAND3x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND3x2_ASAP7_6t_SL 0 0 ; 
  SIZE 4.32 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.612 0.54 4.004 0.612 ; 
        RECT 3.932 0.396 4.004 0.612 ; 
        RECT 3.564 0.396 4.004 0.468 ; 
        RECT 0.612 0.396 0.684 0.612 ; 
        RECT 0.376 0.396 0.684 0.468 ; 
    END 
  END A 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.076 0.252 2.316 0.324 ; 
        RECT 2.076 0.396 2.3 0.468 ; 
        RECT 2.076 0.252 2.148 0.468 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 4.32 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.32 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.684 4.248 0.756 ; 
        RECT 4.176 0.108 4.248 0.756 ; 
        RECT 3.616 0.108 4.248 0.18 ; 
        RECT 0.072 0.108 0.704 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END Y 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 1.24 0.396 3.008 0.468 ; 
      LAYER M1 ; 
        RECT 2.604 0.396 3.008 0.468 ; 
        RECT 2.604 0.252 2.844 0.324 ; 
        RECT 2.604 0.252 2.676 0.468 ; 
        RECT 1.24 0.396 1.716 0.468 ; 
        RECT 1.644 0.252 1.716 0.468 ; 
        RECT 1.476 0.252 1.716 0.324 ; 
      LAYER V1 ; 
        RECT 1.26 0.396 1.332 0.468 ; 
        RECT 2.916 0.396 2.988 0.468 ; 
    END 
  END B 
  OBS 
    LAYER M1 ; 
      RECT 2.968 0.252 3.944 0.324 ; 
      RECT 1.024 0.108 3.296 0.18 ; 
      RECT 0.376 0.252 1.352 0.324 ; 
  END 
END NAND3x2_ASAP7_6t_SL 


MACRO NAND3xp33R_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND3xp33R_ASAP7_6t_SL 0 0 ; 
  SIZE 1.08 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.344 0.54 0.492 0.612 ; 
        RECT 0.344 0.108 0.492 0.256 ; 
        RECT 0.344 0.108 0.416 0.612 ; 
        RECT 0.272 0.4 0.416 0.472 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.54 0.74 0.612 ; 
        RECT 0.588 0.108 0.736 0.256 ; 
        RECT 0.592 0.108 0.664 0.612 ; 
        RECT 0.516 0.384 0.664 0.456 ; 
        RECT 0.588 0.108 0.664 0.456 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.684 1.008 0.756 ; 
        RECT 0.936 0.108 1.008 0.756 ; 
        RECT 0.808 0.108 1.008 0.256 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.08 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.08 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.096 0.684 0.684 0.756 ; 
        RECT 0.096 0.108 0.272 0.256 ; 
        RECT 0.096 0.108 0.168 0.756 ; 
    END 
  END Y 
END NAND3xp33R_ASAP7_6t_SL 


MACRO NAND3xp33_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND3xp33_ASAP7_6t_SL 0 0 ; 
  SIZE 1.08 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.216 0.54 0.38 0.612 ; 
        RECT 0.216 0.252 0.38 0.324 ; 
        RECT 0.216 0.252 0.288 0.612 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.108 0.704 0.256 ; 
        RECT 0.504 0.54 0.652 0.612 ; 
        RECT 0.504 0.108 0.576 0.612 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.604 1.008 0.756 ; 
        RECT 0.936 0.108 1.008 0.756 ; 
        RECT 0.712 0.396 1.008 0.468 ; 
        RECT 0.812 0.108 1.008 0.256 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.08 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.08 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.684 0.704 0.756 ; 
        RECT 0.072 0.108 0.292 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END Y 
END NAND3xp33_ASAP7_6t_SL 


MACRO NAND4xp25R_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND4xp25R_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.968 0.464 1.116 0.612 ; 
        RECT 1.044 0.252 1.116 0.612 ; 
        RECT 0.936 0.252 1.116 0.324 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.648 0.54 0.868 0.612 ; 
        RECT 0.648 0.396 0.868 0.468 ; 
        RECT 0.648 0.108 0.864 0.18 ; 
        RECT 0.648 0.108 0.72 0.612 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.54 0.576 0.612 ; 
        RECT 0.504 0.108 0.576 0.612 ; 
        RECT 0.376 0.108 0.576 0.256 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.076 0.54 0.296 0.612 ; 
        RECT 0.076 0.396 0.296 0.468 ; 
        RECT 0.076 0.108 0.272 0.256 ; 
        RECT 0.076 0.108 0.148 0.612 ; 
    END 
  END D 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.16 0.684 1.26 0.756 ; 
        RECT 1.188 0.108 1.26 0.756 ; 
        RECT 1.024 0.108 1.26 0.18 ; 
    END 
  END Y 
END NAND4xp25R_ASAP7_6t_SL 


MACRO NAND4xp25_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND4xp25_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.9 0.54 1.08 0.612 ; 
        RECT 1.008 0.36 1.08 0.612 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.648 0.108 0.92 0.256 ; 
        RECT 0.648 0.396 0.828 0.468 ; 
        RECT 0.648 0.108 0.72 0.584 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.54 0.576 0.612 ; 
        RECT 0.504 0.108 0.576 0.612 ; 
        RECT 0.36 0.108 0.576 0.28 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.54 0.292 0.612 ; 
        RECT 0.072 0.396 0.292 0.468 ; 
        RECT 0.072 0.108 0.272 0.28 ; 
        RECT 0.072 0.108 0.144 0.612 ; 
    END 
  END D 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.16 0.684 1.224 0.756 ; 
        RECT 1.152 0.108 1.224 0.756 ; 
        RECT 1.024 0.108 1.224 0.18 ; 
    END 
  END Y 
END NAND4xp25_ASAP7_6t_SL 


MACRO NAND4xp75_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND4xp75_ASAP7_6t_SL 0 0 ; 
  SIZE 3.024 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.508 0.54 2.732 0.612 ; 
        RECT 2.66 0.396 2.732 0.612 ; 
        RECT 2.512 0.396 2.732 0.468 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.888 0.54 2.2 0.612 ; 
        RECT 2.124 0.396 2.196 0.612 ; 
        RECT 1.888 0.396 2.196 0.468 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.54 1.336 0.612 ; 
        RECT 1.264 0.396 1.336 0.612 ; 
        RECT 1.024 0.396 1.336 0.468 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.704 0.468 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END D 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.024 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.024 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 2.952 0.756 ; 
        RECT 2.88 0.108 2.952 0.756 ; 
        RECT 2.32 0.108 2.952 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.672 0.252 2.648 0.324 ; 
      RECT 1.024 0.108 2 0.18 ; 
      RECT 0.376 0.252 1.352 0.324 ; 
  END 
END NAND4xp75_ASAP7_6t_SL 


MACRO NAND5xp2R_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND5xp2R_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.18 0.54 0.328 0.612 ; 
        RECT 0.18 0.28 0.252 0.612 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.5 0.108 0.572 0.464 ; 
        RECT 0.376 0.108 0.572 0.256 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.108 0.92 0.256 ; 
        RECT 0.72 0.54 0.868 0.612 ; 
        RECT 0.72 0.108 0.792 0.612 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.02 0.464 1.168 0.612 ; 
        RECT 1.02 0.108 1.168 0.256 ; 
        RECT 0.928 0.392 1.092 0.464 ; 
        RECT 1.02 0.108 1.092 0.612 ; 
    END 
  END D 
  PIN E 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.24 0.608 1.476 0.756 ; 
        RECT 1.404 0.108 1.476 0.756 ; 
        RECT 1.312 0.392 1.476 0.464 ; 
        RECT 1.24 0.108 1.476 0.256 ; 
    END 
  END E 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.036 0.684 1.136 0.756 ; 
        RECT 0.036 0.108 0.272 0.18 ; 
        RECT 0.036 0.108 0.108 0.756 ; 
    END 
  END Y 
END NAND5xp2R_ASAP7_6t_SL 


MACRO NAND5xp2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND5xp2_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.18 0.252 0.476 0.324 ; 
        RECT 0.18 0.54 0.452 0.612 ; 
        RECT 0.18 0.252 0.252 0.612 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.576 0.108 0.648 0.584 ; 
        RECT 0.352 0.396 0.648 0.468 ; 
        RECT 0.396 0.108 0.648 0.18 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.108 0.92 0.272 ; 
        RECT 0.72 0.54 0.908 0.612 ; 
        RECT 0.72 0.108 0.792 0.612 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.008 0.46 1.164 0.612 ; 
        RECT 1.008 0.108 1.156 0.264 ; 
        RECT 0.936 0.392 1.08 0.464 ; 
        RECT 1.008 0.108 1.08 0.612 ; 
    END 
  END D 
  PIN E 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.236 0.604 1.44 0.756 ; 
        RECT 1.368 0.108 1.44 0.756 ; 
        RECT 1.276 0.392 1.44 0.464 ; 
        RECT 1.24 0.108 1.44 0.264 ; 
    END 
  END E 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.036 0.684 1.136 0.756 ; 
        RECT 0.036 0.108 0.272 0.18 ; 
        RECT 0.036 0.108 0.108 0.756 ; 
    END 
  END Y 
END NAND5xp2_ASAP7_6t_SL 


MACRO NOR2x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR2x1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.336 0.468 ; 
        RECT 0.072 0.54 0.292 0.612 ; 
        RECT 0.072 0.108 0.272 0.26 ; 
        RECT 0.072 0.108 0.144 0.612 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.46 0.396 0.92 0.468 ; 
        RECT 0.46 0.54 0.68 0.612 ; 
        RECT 0.46 0.252 0.68 0.324 ; 
        RECT 0.46 0.252 0.532 0.612 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.54 1.244 0.612 ; 
        RECT 1.172 0.108 1.244 0.612 ; 
        RECT 0.376 0.108 1.244 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.684 1.136 0.756 ; 
  END 
END NOR2x1_ASAP7_6t_SL 


MACRO NOR2x2R_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR2x2R_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.468 0.468 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.612 0.396 1.12 0.468 ; 
        RECT 0.532 0.54 0.684 0.612 ; 
        RECT 0.612 0.252 0.684 0.612 ; 
        RECT 0.536 0.252 0.684 0.324 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.044 0.684 1.656 0.756 ; 
        RECT 1.584 0.108 1.656 0.756 ; 
        RECT 0.376 0.108 1.656 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.808 0.54 1.352 0.612 ; 
      RECT 0.376 0.684 0.92 0.756 ; 
  END 
END NOR2x2R_ASAP7_6t_SL 


MACRO NOR2x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR2x2_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.968 0.396 1.188 0.468 ; 
        RECT 1.116 0.252 1.188 0.468 ; 
        RECT 0.968 0.252 1.188 0.324 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.288 0.396 1.872 0.468 ; 
        RECT 1.8 0.252 1.872 0.468 ; 
        RECT 1.652 0.252 1.872 0.324 ; 
        RECT 0.728 0.54 1.36 0.612 ; 
        RECT 1.288 0.396 1.36 0.612 ; 
        RECT 0.728 0.396 0.8 0.612 ; 
        RECT 0.288 0.396 0.8 0.468 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.672 0.54 2.088 0.612 ; 
        RECT 2.016 0.108 2.088 0.612 ; 
        RECT 0.072 0.108 2.088 0.18 ; 
        RECT 0.072 0.54 0.488 0.612 ; 
        RECT 0.072 0.108 0.144 0.612 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.684 2 0.756 ; 
  END 
END NOR2x2_ASAP7_6t_SL 


MACRO NOR2xp5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR2xp5_ASAP7_6t_SL 0 0 ; 
  SIZE 0.864 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.068 0.412 0.308 0.484 ; 
        RECT 0.068 0.608 0.272 0.756 ; 
        RECT 0.068 0.108 0.272 0.18 ; 
        RECT 0.068 0.108 0.14 0.756 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.416 0.396 0.596 0.468 ; 
        RECT 0.344 0.608 0.492 0.756 ; 
        RECT 0.416 0.396 0.492 0.756 ; 
        RECT 0.416 0.252 0.488 0.756 ; 
        RECT 0.34 0.252 0.488 0.324 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 0.864 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.864 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.684 0.792 0.756 ; 
        RECT 0.72 0.108 0.792 0.756 ; 
        RECT 0.396 0.108 0.792 0.18 ; 
    END 
  END Y 
END NOR2xp5_ASAP7_6t_SL 


MACRO NOR3x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR3x1_ASAP7_6t_SL 0 0 ; 
  SIZE 2.376 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.396 1.872 0.468 ; 
        RECT 1.8 0.252 1.872 0.468 ; 
        RECT 1.584 0.252 1.872 0.324 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.532 0.396 1.352 0.468 ; 
        RECT 0.532 0.54 0.9 0.612 ; 
        RECT 0.532 0.108 0.708 0.284 ; 
        RECT 0.532 0.108 0.604 0.612 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.316 0.468 ; 
        RECT 0.072 0.108 0.292 0.18 ; 
        RECT 0.072 0.588 0.272 0.756 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.376 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.672 0.684 2.304 0.756 ; 
        RECT 2.232 0.108 2.304 0.756 ; 
        RECT 0.808 0.108 2.304 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.024 0.54 2 0.612 ; 
      RECT 0.376 0.684 1.352 0.756 ; 
  END 
END NOR3x1_ASAP7_6t_SL 


MACRO NOR3x1f_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR3x1f_ASAP7_6t_SL 0 0 ; 
  SIZE 1.08 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.344 0.608 0.492 0.756 ; 
        RECT 0.344 0.252 0.492 0.324 ; 
        RECT 0.344 0.252 0.416 0.756 ; 
        RECT 0.252 0.396 0.416 0.468 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.252 0.74 0.324 ; 
        RECT 0.588 0.556 0.736 0.756 ; 
        RECT 0.588 0.408 0.664 0.756 ; 
        RECT 0.592 0.252 0.664 0.756 ; 
        RECT 0.516 0.408 0.664 0.48 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.556 1.008 0.756 ; 
        RECT 0.936 0.108 1.008 0.756 ; 
        RECT 0.808 0.108 1.008 0.18 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.08 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.08 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 0.684 0.18 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END Y 
END NOR3x1f_ASAP7_6t_SL 


MACRO NOR3x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR3x2_ASAP7_6t_SL 0 0 ; 
  SIZE 4.32 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 3.784 0.396 4.004 0.468 ; 
        RECT 3.932 0.252 4.004 0.468 ; 
        RECT 0.612 0.252 4.004 0.324 ; 
        RECT 0.376 0.396 0.684 0.468 ; 
        RECT 0.612 0.252 0.684 0.468 ; 
    END 
  END A 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.076 0.54 2.316 0.612 ; 
        RECT 2.076 0.396 2.3 0.468 ; 
        RECT 2.076 0.396 2.148 0.612 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 4.32 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.32 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 3.52 0.684 4.248 0.756 ; 
        RECT 4.176 0.108 4.248 0.756 ; 
        RECT 0.072 0.108 4.248 0.18 ; 
        RECT 0.072 0.684 0.704 0.756 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END Y 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 1.24 0.396 3.008 0.468 ; 
      LAYER M1 ; 
        RECT 2.604 0.396 3.008 0.468 ; 
        RECT 2.604 0.54 2.844 0.612 ; 
        RECT 2.604 0.396 2.676 0.612 ; 
        RECT 1.476 0.54 1.716 0.612 ; 
        RECT 1.644 0.396 1.716 0.612 ; 
        RECT 1.24 0.396 1.716 0.468 ; 
      LAYER V1 ; 
        RECT 1.26 0.396 1.332 0.468 ; 
        RECT 2.916 0.396 2.988 0.468 ; 
    END 
  END B 
  OBS 
    LAYER M1 ; 
      RECT 2.968 0.54 3.944 0.612 ; 
      RECT 1.024 0.684 3.296 0.756 ; 
      RECT 0.376 0.54 1.352 0.612 ; 
  END 
END NOR3x2_ASAP7_6t_SL 


MACRO NOR3xp33_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR3xp33_ASAP7_6t_SL 0 0 ; 
  SIZE 1.08 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.344 0.608 0.492 0.756 ; 
        RECT 0.344 0.252 0.492 0.324 ; 
        RECT 0.344 0.252 0.416 0.756 ; 
        RECT 0.252 0.396 0.416 0.468 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.252 0.74 0.324 ; 
        RECT 0.588 0.556 0.736 0.756 ; 
        RECT 0.588 0.408 0.664 0.756 ; 
        RECT 0.592 0.252 0.664 0.756 ; 
        RECT 0.516 0.408 0.664 0.48 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.556 1.008 0.756 ; 
        RECT 0.936 0.108 1.008 0.756 ; 
        RECT 0.808 0.108 1.008 0.18 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.08 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.08 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 0.684 0.18 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END Y 
END NOR3xp33_ASAP7_6t_SL 


MACRO NOR4x3f_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR4x3f_ASAP7_6t_SL 0 0 ; 
  SIZE 3.024 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.3 0.396 2.58 0.468 ; 
        RECT 2.508 0.252 2.58 0.468 ; 
        RECT 1.948 0.252 2.58 0.324 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.412 0.396 2.004 0.468 ; 
        RECT 1.412 0.252 1.584 0.612 ; 
        RECT 1.056 0.252 1.584 0.324 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.612 0.396 1.16 0.468 ; 
        RECT 0.372 0.54 0.684 0.612 ; 
        RECT 0.612 0.252 0.684 0.612 ; 
        RECT 0.376 0.252 0.684 0.324 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.468 0.468 ; 
        RECT 0.072 0.108 0.272 0.26 ; 
        RECT 0.072 0.596 0.268 0.756 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END D 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.024 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.024 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.32 0.684 2.952 0.756 ; 
        RECT 2.88 0.108 2.952 0.756 ; 
        RECT 0.376 0.108 2.952 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.368 0.684 0.864 0.756 ; 
      RECT 0.792 0.54 0.864 0.756 ; 
      RECT 0.792 0.54 1.312 0.612 ; 
      RECT 1.712 0.54 2.664 0.612 ; 
      RECT 1 0.684 2 0.756 ; 
  END 
END NOR4x3f_ASAP7_6t_SL 


MACRO NOR4xp25_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR4xp25_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.008 0.252 1.08 0.504 ; 
        RECT 0.9 0.252 1.08 0.324 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.648 0.608 0.92 0.756 ; 
        RECT 0.648 0.396 0.828 0.468 ; 
        RECT 0.648 0.352 0.72 0.756 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.36 0.584 0.576 0.756 ; 
        RECT 0.504 0.252 0.576 0.756 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.292 0.468 ; 
        RECT 0.072 0.252 0.292 0.324 ; 
        RECT 0.072 0.584 0.272 0.756 ; 
        RECT 0.072 0.252 0.144 0.756 ; 
    END 
  END D 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.684 1.224 0.756 ; 
        RECT 1.152 0.108 1.224 0.756 ; 
        RECT 0.16 0.108 1.224 0.18 ; 
    END 
  END Y 
END NOR4xp25_ASAP7_6t_SL 


MACRO NOR5x1f_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR5x1f_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.684 0.296 0.756 ; 
        RECT 0.072 0.172 0.144 0.756 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.42 0.684 0.576 0.756 ; 
        RECT 0.504 0.252 0.576 0.756 ; 
        RECT 0.392 0.252 0.576 0.324 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.648 0.6 0.868 0.756 ; 
        RECT 0.648 0.252 0.868 0.408 ; 
        RECT 0.72 0.252 0.792 0.756 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.94 0.252 1.248 0.324 ; 
        RECT 0.94 0.684 1.172 0.756 ; 
        RECT 0.94 0.252 1.012 0.756 ; 
    END 
  END D 
  PIN E 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.296 0.684 1.444 0.756 ; 
        RECT 1.372 0.108 1.444 0.756 ; 
        RECT 1.296 0.108 1.444 0.18 ; 
    END 
  END E 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.22 0.108 1.14 0.18 ; 
        RECT 0.22 0.54 0.384 0.612 ; 
        RECT 0.22 0.108 0.292 0.612 ; 
    END 
  END Y 
END NOR5x1f_ASAP7_6t_SL 


MACRO NOR5xp2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR5xp2_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.18 0.54 0.476 0.612 ; 
        RECT 0.18 0.252 0.452 0.324 ; 
        RECT 0.18 0.252 0.252 0.612 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.684 0.648 0.756 ; 
        RECT 0.576 0.28 0.648 0.756 ; 
        RECT 0.352 0.396 0.648 0.468 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.592 0.92 0.756 ; 
        RECT 0.72 0.252 0.908 0.324 ; 
        RECT 0.72 0.252 0.792 0.756 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.008 0.252 1.164 0.404 ; 
        RECT 1.008 0.6 1.156 0.756 ; 
        RECT 1.008 0.252 1.08 0.756 ; 
        RECT 0.936 0.4 1.08 0.472 ; 
    END 
  END D 
  PIN E 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.24 0.6 1.44 0.756 ; 
        RECT 1.368 0.108 1.44 0.756 ; 
        RECT 1.276 0.4 1.44 0.472 ; 
        RECT 1.236 0.108 1.44 0.26 ; 
    END 
  END E 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.036 0.108 1.136 0.18 ; 
        RECT 0.036 0.684 0.272 0.756 ; 
        RECT 0.036 0.108 0.108 0.756 ; 
    END 
  END Y 
END NOR5xp2_ASAP7_6t_SL 


MACRO O2A1O1A1Ixp33_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN O2A1O1A1Ixp33_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.684 0.22 0.756 ; 
        RECT 0.072 0.252 0.22 0.324 ; 
        RECT 0.072 0.252 0.144 0.756 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.42 0.396 0.576 0.468 ; 
        RECT 0.344 0.54 0.492 0.612 ; 
        RECT 0.42 0.256 0.492 0.612 ; 
        RECT 0.344 0.256 0.492 0.328 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.54 0.872 0.612 ; 
        RECT 0.72 0.252 0.872 0.324 ; 
        RECT 0.72 0.252 0.792 0.612 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.148 0.54 1.3 0.612 ; 
        RECT 1.148 0.252 1.3 0.324 ; 
        RECT 1.148 0.252 1.22 0.612 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.504 0.54 1.656 0.612 ; 
        RECT 1.584 0.256 1.656 0.612 ; 
        RECT 1.504 0.256 1.656 0.328 ; 
    END 
  END D 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.044 0.684 1.872 0.756 ; 
        RECT 1.8 0.108 1.872 0.756 ; 
        RECT 1.692 0.108 1.872 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.828 0.108 1.548 0.18 ; 
      RECT 0.396 0.684 0.9 0.756 ; 
      RECT 0.16 0.108 0.684 0.18 ; 
  END 
END O2A1O1A1Ixp33_ASAP7_6t_SL 


MACRO O2A1O1Ixp33_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN O2A1O1Ixp33_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.684 0.272 0.756 ; 
        RECT 0.072 0.252 0.224 0.4 ; 
        RECT 0.072 0.252 0.144 0.756 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.4 0.396 0.568 0.468 ; 
        RECT 0.324 0.54 0.472 0.612 ; 
        RECT 0.4 0.252 0.472 0.612 ; 
        RECT 0.324 0.252 0.472 0.4 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.616 0.54 0.78 0.612 ; 
        RECT 0.708 0.252 0.78 0.612 ; 
        RECT 0.616 0.252 0.78 0.324 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.996 0.252 1.068 0.544 ; 
        RECT 0.86 0.464 1.008 0.612 ; 
        RECT 0.88 0.252 1.068 0.324 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.044 0.684 1.26 0.756 ; 
        RECT 1.188 0.108 1.26 0.756 ; 
        RECT 0.828 0.108 1.26 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.396 0.684 0.9 0.756 ; 
      RECT 0.16 0.108 0.684 0.18 ; 
  END 
END O2A1O1Ixp33_ASAP7_6t_SL 


MACRO O2A1O1Ixp5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN O2A1O1Ixp5_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.928 0.252 1 0.416 ; 
        RECT 0.072 0.252 1 0.324 ; 
        RECT 0.072 0.108 0.468 0.18 ; 
        RECT 0.072 0.684 0.272 0.756 ; 
        RECT 0.072 0.108 0.148 0.324 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.34 0.396 0.704 0.468 ; 
        RECT 0.34 0.396 0.488 0.612 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.184 0.252 1.376 0.324 ; 
        RECT 1.164 0.256 1.236 0.488 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.324 0.54 1.52 0.612 ; 
        RECT 1.448 0.376 1.52 0.612 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.592 0.108 1.664 0.628 ; 
        RECT 1.26 0.108 1.664 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.024 0.684 1.332 0.756 ; 
      RECT 1.024 0.54 1.096 0.756 ; 
      RECT 0.612 0.54 1.096 0.612 ; 
      RECT 0.592 0.108 1.136 0.18 ; 
      RECT 0.396 0.684 0.9 0.756 ; 
  END 
END O2A1O1Ixp5_ASAP7_6t_SL 


MACRO OA211x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA211x1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.456 0.54 0.612 0.612 ; 
        RECT 0.516 0.384 0.588 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.064 0.684 0.212 0.756 ; 
        RECT 0.14 0.252 0.212 0.756 ; 
        RECT 0.064 0.252 0.212 0.324 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.016 0.108 1.136 0.256 ; 
        RECT 0.936 0.396 1.088 0.468 ; 
        RECT 1.016 0.108 1.088 0.468 ; 
        RECT 0.936 0.108 1.136 0.18 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.712 0.252 0.892 0.324 ; 
        RECT 0.712 0.54 0.864 0.612 ; 
        RECT 0.712 0.252 0.784 0.612 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.196 0.684 1.476 0.756 ; 
        RECT 1.404 0.108 1.476 0.756 ; 
        RECT 1.24 0.108 1.476 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.284 0.684 1.072 0.756 ; 
      RECT 1 0.54 1.072 0.756 ; 
      RECT 0.284 0.252 0.356 0.756 ; 
      RECT 1 0.54 1.232 0.612 ; 
      RECT 1.16 0.372 1.232 0.612 ; 
      RECT 1.16 0.396 1.304 0.468 ; 
      RECT 0.284 0.252 0.432 0.324 ; 
      RECT 0.16 0.108 0.756 0.18 ; 
  END 
END OA211x1_ASAP7_6t_SL 


MACRO OA211x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA211x2_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.456 0.54 0.612 0.612 ; 
        RECT 0.516 0.36 0.588 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.064 0.684 0.212 0.756 ; 
        RECT 0.14 0.252 0.212 0.756 ; 
        RECT 0.064 0.252 0.212 0.324 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.016 0.108 1.24 0.304 ; 
        RECT 0.936 0.396 1.088 0.468 ; 
        RECT 1.016 0.108 1.088 0.468 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.712 0.54 1.06 0.612 ; 
        RECT 0.712 0.252 0.892 0.324 ; 
        RECT 0.712 0.252 0.784 0.612 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.312 0.684 1.648 0.756 ; 
        RECT 1.576 0.108 1.648 0.756 ; 
        RECT 1.312 0.108 1.648 0.18 ; 
        RECT 1.312 0.588 1.384 0.756 ; 
        RECT 1.312 0.108 1.384 0.272 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.284 0.684 1.236 0.756 ; 
      RECT 1.164 0.396 1.236 0.756 ; 
      RECT 0.284 0.252 0.356 0.756 ; 
      RECT 1.164 0.396 1.384 0.468 ; 
      RECT 0.284 0.252 0.432 0.324 ; 
      RECT 0.14 0.108 0.772 0.18 ; 
  END 
END OA211x2_ASAP7_6t_SL 


MACRO OA21x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21x1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.068 0.684 0.272 0.756 ; 
        RECT 0.068 0.38 0.14 0.756 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.532 0.54 0.68 0.612 ; 
        RECT 0.532 0.252 0.68 0.324 ; 
        RECT 0.532 0.252 0.604 0.612 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.804 0.464 0.952 0.612 ; 
        RECT 0.804 0.108 0.952 0.256 ; 
        RECT 0.732 0.396 0.876 0.468 ; 
        RECT 0.804 0.108 0.876 0.612 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.188 0.108 1.26 0.672 ; 
        RECT 1.024 0.108 1.26 0.256 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.372 0.684 1.116 0.756 ; 
      RECT 1.044 0.376 1.116 0.756 ; 
      RECT 0.372 0.532 0.444 0.756 ; 
      RECT 0.284 0.532 0.444 0.604 ; 
      RECT 0.284 0.252 0.356 0.604 ; 
      RECT 0.284 0.252 0.432 0.324 ; 
      RECT 0.16 0.108 0.704 0.18 ; 
  END 
END OA21x1_ASAP7_6t_SL 


MACRO OA21x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21x2_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.064 0.684 0.272 0.756 ; 
        RECT 0.064 0.38 0.136 0.756 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.532 0.54 0.68 0.612 ; 
        RECT 0.532 0.252 0.68 0.324 ; 
        RECT 0.532 0.252 0.604 0.612 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.804 0.464 0.952 0.612 ; 
        RECT 0.804 0.108 0.952 0.18 ; 
        RECT 0.728 0.396 0.876 0.468 ; 
        RECT 0.804 0.108 0.876 0.612 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.172 0.108 1.404 0.18 ; 
        RECT 1.052 0.54 1.244 0.612 ; 
        RECT 1.172 0.108 1.244 0.612 ; 
        RECT 1.032 0.252 1.244 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.372 0.684 1.436 0.756 ; 
      RECT 1.364 0.376 1.436 0.756 ; 
      RECT 0.372 0.532 0.444 0.756 ; 
      RECT 0.284 0.532 0.444 0.604 ; 
      RECT 0.284 0.252 0.36 0.604 ; 
      RECT 0.284 0.252 0.432 0.324 ; 
      RECT 0.16 0.108 0.684 0.18 ; 
  END 
END OA21x2_ASAP7_6t_SL 


MACRO OA221x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA221x1_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.32 0.396 0.576 0.468 ; 
        RECT 0.32 0.684 0.468 0.756 ; 
        RECT 0.32 0.252 0.468 0.468 ; 
        RECT 0.32 0.252 0.392 0.756 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.684 0.22 0.756 ; 
        RECT 0.072 0.252 0.22 0.324 ; 
        RECT 0.072 0.252 0.144 0.756 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.48 0.108 1.764 0.26 ; 
        RECT 1.444 0.54 1.612 0.612 ; 
        RECT 1.48 0.108 1.552 0.612 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.856 0.54 1.172 0.612 ; 
        RECT 0.856 0.396 1.172 0.468 ; 
        RECT 0.856 0.284 0.928 0.612 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.536 0.54 0.784 0.612 ; 
        RECT 0.712 0.252 0.784 0.612 ; 
        RECT 0.612 0.252 0.784 0.324 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.888 0.684 2.064 0.756 ; 
        RECT 1.992 0.108 2.064 0.756 ; 
        RECT 1.888 0.108 2.064 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.592 0.684 1.788 0.756 ; 
      RECT 1.716 0.396 1.788 0.756 ; 
      RECT 1.272 0.252 1.344 0.756 ; 
      RECT 1.716 0.396 1.892 0.468 ; 
      RECT 1.064 0.252 1.344 0.324 ; 
      RECT 0.828 0.108 1.332 0.18 ; 
      RECT 0.16 0.108 0.684 0.18 ; 
  END 
END OA221x1_ASAP7_6t_SL 


MACRO OA221x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA221x2_ASAP7_6t_SL 0 0 ; 
  SIZE 2.376 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.32 0.396 0.576 0.468 ; 
        RECT 0.32 0.684 0.468 0.756 ; 
        RECT 0.32 0.252 0.468 0.468 ; 
        RECT 0.32 0.252 0.392 0.756 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.684 0.22 0.756 ; 
        RECT 0.072 0.252 0.22 0.324 ; 
        RECT 0.072 0.252 0.144 0.756 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.48 0.108 1.764 0.26 ; 
        RECT 1.444 0.54 1.612 0.612 ; 
        RECT 1.48 0.108 1.552 0.612 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.856 0.54 1.172 0.612 ; 
        RECT 0.856 0.396 1.172 0.468 ; 
        RECT 0.856 0.284 0.928 0.612 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.536 0.54 0.784 0.612 ; 
        RECT 0.712 0.252 0.784 0.612 ; 
        RECT 0.612 0.252 0.784 0.324 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.376 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.888 0.684 2.204 0.756 ; 
        RECT 2.124 0.108 2.204 0.756 ; 
        RECT 1.888 0.108 2.204 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.592 0.684 1.788 0.756 ; 
      RECT 1.716 0.396 1.788 0.756 ; 
      RECT 1.272 0.252 1.344 0.756 ; 
      RECT 1.716 0.396 1.892 0.468 ; 
      RECT 1.064 0.252 1.344 0.324 ; 
      RECT 0.828 0.108 1.332 0.18 ; 
      RECT 0.16 0.108 0.684 0.18 ; 
  END 
END OA221x2_ASAP7_6t_SL 


MACRO OA222x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA222x1_ASAP7_6t_SL 0 0 ; 
  SIZE 2.376 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.096 0.684 0.276 0.756 ; 
        RECT 0.204 0.252 0.276 0.756 ; 
        RECT 0.096 0.252 0.276 0.324 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.496 0.54 0.668 0.612 ; 
        RECT 0.496 0.252 0.668 0.324 ; 
        RECT 0.496 0.252 0.568 0.612 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.132 0.54 1.352 0.612 ; 
        RECT 1.28 0.396 1.352 0.612 ; 
        RECT 1.132 0.396 1.352 0.468 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.792 0.54 1.012 0.612 ; 
        RECT 0.94 0.396 1.012 0.612 ; 
        RECT 0.72 0.396 1.012 0.468 ; 
    END 
  END B2 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.432 0.54 1.656 0.612 ; 
        RECT 1.432 0.396 1.656 0.468 ; 
        RECT 1.432 0.396 1.504 0.612 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.76 0.464 1.92 0.612 ; 
        RECT 1.8 0.252 1.872 0.612 ; 
        RECT 1.644 0.252 1.872 0.324 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.376 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.192 0.608 2.34 0.756 ; 
        RECT 2.192 0.108 2.34 0.256 ; 
        RECT 2.192 0.108 2.264 0.756 ; 
        RECT 2.1 0.108 2.34 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.348 0.684 2.092 0.756 ; 
      RECT 2.02 0.376 2.092 0.756 ; 
      RECT 0.348 0.232 0.42 0.756 ; 
      RECT 0.844 0.252 1.44 0.324 ; 
      RECT 1.368 0.108 1.44 0.324 ; 
      RECT 1.368 0.108 1.784 0.18 ; 
      RECT 1.024 0.108 1.236 0.18 ; 
      RECT 0.592 0.108 0.74 0.18 ; 
      RECT 0.072 0.108 0.272 0.18 ; 
    LAYER M2 ; 
      RECT 0.16 0.108 1.148 0.18 ; 
    LAYER V1 ; 
      RECT 1.044 0.108 1.116 0.18 ; 
      RECT 0.612 0.108 0.684 0.18 ; 
      RECT 0.18 0.108 0.252 0.18 ; 
  END 
END OA222x1_ASAP7_6t_SL 


MACRO OA222x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA222x2_ASAP7_6t_SL 0 0 ; 
  SIZE 2.592 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.064 0.396 0.28 0.468 ; 
        RECT 0.208 0.304 0.28 0.468 ; 
        RECT 0.064 0.608 0.272 0.756 ; 
        RECT 0.064 0.396 0.136 0.756 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.496 0.54 0.668 0.612 ; 
        RECT 0.496 0.252 0.648 0.324 ; 
        RECT 0.496 0.252 0.568 0.612 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.132 0.54 1.352 0.612 ; 
        RECT 1.28 0.396 1.352 0.612 ; 
        RECT 1.132 0.396 1.352 0.468 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.8 0.396 1.012 0.604 ; 
        RECT 0.728 0.396 1.012 0.468 ; 
    END 
  END B2 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.432 0.54 1.656 0.612 ; 
        RECT 1.432 0.396 1.656 0.468 ; 
        RECT 1.432 0.396 1.504 0.612 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.76 0.464 1.928 0.612 ; 
        RECT 1.8 0.252 1.872 0.612 ; 
        RECT 1.644 0.252 1.872 0.324 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.592 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.176 0.684 2.52 0.756 ; 
        RECT 2.448 0.108 2.52 0.756 ; 
        RECT 2.104 0.108 2.52 0.18 ; 
        RECT 2.176 0.568 2.248 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.352 0.684 2.104 0.756 ; 
      RECT 2.032 0.396 2.104 0.756 ; 
      RECT 0.352 0.184 0.424 0.756 ; 
      RECT 0.844 0.252 1.44 0.324 ; 
      RECT 1.368 0.108 1.44 0.324 ; 
      RECT 1.368 0.108 1.872 0.18 ; 
      RECT 0.072 0.108 0.144 0.256 ; 
      RECT 0.072 0.108 0.26 0.18 ; 
      RECT 1.024 0.108 1.236 0.18 ; 
      RECT 0.592 0.108 0.74 0.18 ; 
    LAYER M2 ; 
      RECT 0.08 0.108 1.148 0.18 ; 
    LAYER V1 ; 
      RECT 1.044 0.108 1.116 0.18 ; 
      RECT 0.612 0.108 0.684 0.18 ; 
      RECT 0.18 0.108 0.252 0.18 ; 
  END 
END OA222x2_ASAP7_6t_SL 


MACRO OA22x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA22x1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.124 0.684 0.272 0.756 ; 
        RECT 0.2 0.252 0.272 0.756 ; 
        RECT 0.124 0.252 0.272 0.324 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.42 0.4 0.564 0.472 ; 
        RECT 0.344 0.608 0.492 0.756 ; 
        RECT 0.42 0.252 0.492 0.756 ; 
        RECT 0.344 0.252 0.492 0.4 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.236 0.54 1.384 0.612 ; 
        RECT 1.236 0.108 1.384 0.18 ; 
        RECT 1.236 0.108 1.308 0.612 ; 
        RECT 1.164 0.396 1.308 0.468 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.604 0.768 0.756 ; 
        RECT 0.696 0.252 0.768 0.756 ; 
        RECT 0.62 0.252 0.768 0.324 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.672 0.684 1.832 0.756 ; 
        RECT 1.76 0.108 1.832 0.756 ; 
        RECT 1.672 0.108 1.832 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.94 0.684 1.572 0.756 ; 
      RECT 1.5 0.396 1.572 0.756 ; 
      RECT 0.94 0.252 1.016 0.756 ; 
      RECT 0.868 0.576 1.016 0.648 ; 
      RECT 1.5 0.396 1.66 0.468 ; 
      RECT 0.868 0.252 1.016 0.324 ; 
      RECT 0.16 0.108 1.136 0.18 ; 
  END 
END OA22x1_ASAP7_6t_SL 


MACRO OA22x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA22x2_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.944 0.684 2.092 0.756 ; 
        RECT 2.02 0.252 2.092 0.756 ; 
        RECT 1.944 0.252 2.092 0.324 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.696 0.608 1.844 0.756 ; 
        RECT 1.772 0.252 1.844 0.756 ; 
        RECT 1.596 0.252 1.844 0.324 ; 
        RECT 1.596 0.252 1.668 0.468 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.648 0.396 1 0.468 ; 
        RECT 0.648 0.108 0.8 0.612 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.448 0.604 1.596 0.756 ; 
        RECT 1.448 0.396 1.52 0.756 ; 
        RECT 1.356 0.396 1.52 0.468 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.092 0.68 0.432 0.756 ; 
        RECT 0.36 0.108 0.432 0.756 ; 
        RECT 0.092 0.108 0.432 0.184 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.504 0.684 1.172 0.756 ; 
      RECT 1.1 0.252 1.172 0.756 ; 
      RECT 1.1 0.612 1.32 0.684 ; 
      RECT 0.504 0.356 0.576 0.756 ; 
      RECT 1.1 0.252 1.32 0.324 ; 
      RECT 1 0.108 2.024 0.18 ; 
  END 
END OA22x2_ASAP7_6t_SL 


MACRO OA311x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA311x1_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.54 0.868 0.612 ; 
        RECT 0.72 0.376 0.792 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.576 0.756 ; 
        RECT 0.504 0.252 0.576 0.756 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.404 0.372 0.476 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A3 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.252 1.008 0.488 ; 
        RECT 0.86 0.252 1.008 0.324 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.076 0.54 1.224 0.612 ; 
        RECT 1.152 0.28 1.224 0.612 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.888 0.684 2.084 0.756 ; 
        RECT 2.012 0.108 2.084 0.756 ; 
        RECT 1.888 0.108 2.084 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.792 0.684 1.44 0.756 ; 
      RECT 1.368 0.108 1.44 0.756 ; 
      RECT 1.368 0.396 1.892 0.468 ; 
      RECT 1.24 0.108 1.44 0.18 ; 
      RECT 0.376 0.108 0.936 0.18 ; 
  END 
END OA311x1_ASAP7_6t_SL 


MACRO OA311x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA311x2_ASAP7_6t_SL 0 0 ; 
  SIZE 2.376 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.54 0.868 0.612 ; 
        RECT 0.72 0.376 0.792 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.576 0.756 ; 
        RECT 0.504 0.252 0.576 0.756 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.404 0.372 0.476 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A3 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.252 1.008 0.488 ; 
        RECT 0.86 0.252 1.008 0.324 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.076 0.54 1.224 0.612 ; 
        RECT 1.152 0.28 1.224 0.612 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.376 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.888 0.684 2.3 0.756 ; 
        RECT 2.228 0.108 2.3 0.756 ; 
        RECT 1.888 0.108 2.3 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.792 0.684 1.44 0.756 ; 
      RECT 1.368 0.108 1.44 0.756 ; 
      RECT 1.368 0.396 1.892 0.468 ; 
      RECT 1.24 0.108 1.44 0.18 ; 
      RECT 0.376 0.108 0.936 0.18 ; 
  END 
END OA311x2_ASAP7_6t_SL 


MACRO OA31x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA31x1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.46 0.464 0.612 0.612 ; 
        RECT 0.492 0.252 0.564 0.612 ; 
        RECT 0.392 0.252 0.564 0.324 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.712 0.54 0.888 0.612 ; 
        RECT 0.696 0.252 0.844 0.324 ; 
        RECT 0.712 0.252 0.784 0.612 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.02 0.108 1.168 0.256 ; 
        RECT 0.924 0.396 1.092 0.468 ; 
        RECT 1.02 0.108 1.092 0.468 ; 
    END 
  END A3 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.068 0.684 0.216 0.756 ; 
        RECT 0.068 0.232 0.14 0.756 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.22 0.684 1.44 0.756 ; 
        RECT 1.368 0.108 1.44 0.756 ; 
        RECT 1.292 0.108 1.44 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.316 0.684 1.096 0.756 ; 
      RECT 1.024 0.54 1.096 0.756 ; 
      RECT 0.316 0.496 0.388 0.756 ; 
      RECT 1.024 0.54 1.296 0.612 ; 
      RECT 1.224 0.376 1.296 0.612 ; 
      RECT 0.22 0.496 0.388 0.568 ; 
      RECT 0.22 0.232 0.292 0.568 ; 
      RECT 0.376 0.108 0.92 0.18 ; 
  END 
END OA31x1_ASAP7_6t_SL 


MACRO OA31x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA31x2_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.46 0.464 0.608 0.612 ; 
        RECT 0.492 0.252 0.564 0.612 ; 
        RECT 0.392 0.252 0.564 0.324 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.712 0.54 0.9 0.612 ; 
        RECT 0.68 0.252 0.828 0.4 ; 
        RECT 0.712 0.252 0.784 0.612 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.016 0.108 1.236 0.304 ; 
        RECT 0.936 0.396 1.088 0.468 ; 
        RECT 1.016 0.108 1.088 0.468 ; 
    END 
  END A3 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.068 0.684 0.216 0.756 ; 
        RECT 0.068 0.144 0.14 0.756 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.312 0.684 1.648 0.756 ; 
        RECT 1.576 0.108 1.648 0.756 ; 
        RECT 1.312 0.108 1.648 0.18 ; 
        RECT 1.312 0.588 1.384 0.756 ; 
        RECT 1.312 0.108 1.384 0.272 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.316 0.684 1.232 0.756 ; 
      RECT 1.16 0.396 1.232 0.756 ; 
      RECT 0.316 0.496 0.388 0.756 ; 
      RECT 0.22 0.496 0.388 0.604 ; 
      RECT 0.22 0.232 0.292 0.604 ; 
      RECT 1.16 0.396 1.38 0.468 ; 
      RECT 0.376 0.108 0.9 0.18 ; 
  END 
END OA31x2_ASAP7_6t_SL 


MACRO OA321x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA321x1_ASAP7_6t_SL 0 0 ; 
  SIZE 2.376 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.376 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.376 0.792 0.584 ; 
      LAYER M2 ; 
        RECT 0.632 0.396 0.888 0.468 ; 
      LAYER V1 ; 
        RECT 0.72 0.396 0.792 0.468 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.576 0.756 ; 
        RECT 0.504 0.252 0.576 0.756 ; 
        RECT 0.392 0.252 0.576 0.324 ; 
      LAYER M2 ; 
        RECT 0.388 0.54 0.652 0.612 ; 
      LAYER V1 ; 
        RECT 0.504 0.54 0.576 0.612 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
      LAYER M2 ; 
        RECT 0.072 0.396 0.328 0.468 ; 
      LAYER V1 ; 
        RECT 0.072 0.396 0.144 0.468 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.108 0.684 1.268 0.756 ; 
        RECT 1.152 0.396 1.224 0.756 ; 
      LAYER M2 ; 
        RECT 1.028 0.54 1.344 0.612 ; 
      LAYER V1 ; 
        RECT 1.152 0.54 1.224 0.612 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.54 1.588 0.612 ; 
        RECT 1.368 0.396 1.588 0.468 ; 
        RECT 1.368 0.396 1.44 0.612 ; 
      LAYER M2 ; 
        RECT 1.312 0.396 1.612 0.468 ; 
      LAYER V1 ; 
        RECT 1.388 0.396 1.46 0.468 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.252 1.084 0.324 ; 
        RECT 0.936 0.252 1.008 0.584 ; 
      LAYER M2 ; 
        RECT 0.848 0.252 1.112 0.324 ; 
      LAYER V1 ; 
        RECT 0.956 0.252 1.028 0.324 ; 
    END 
  END C 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.104 0.684 2.3 0.756 ; 
        RECT 2.228 0.108 2.3 0.756 ; 
        RECT 2.104 0.108 2.3 0.18 ; 
      LAYER M2 ; 
        RECT 1.488 0.108 2.3 0.18 ; 
      LAYER V1 ; 
        RECT 2.124 0.108 2.196 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.4 0.684 1.784 0.756 ; 
      RECT 1.712 0.252 1.784 0.756 ; 
      RECT 1.712 0.396 2.108 0.468 ; 
      RECT 1.26 0.252 1.784 0.324 ; 
      RECT 1.024 0.108 1.584 0.18 ; 
      RECT 0.792 0.684 0.952 0.756 ; 
      RECT 0.376 0.108 0.9 0.18 ; 
    LAYER M2 ; 
      RECT 0.828 0.684 1.764 0.756 ; 
    LAYER V1 ; 
      RECT 1.692 0.684 1.764 0.756 ; 
      RECT 0.828 0.684 0.9 0.756 ; 
  END 
END OA321x1_ASAP7_6t_SL 


MACRO OA321x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA321x2_ASAP7_6t_SL 0 0 ; 
  SIZE 2.592 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.592 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.376 0.792 0.584 ; 
      LAYER M2 ; 
        RECT 0.632 0.396 0.888 0.468 ; 
      LAYER V1 ; 
        RECT 0.72 0.396 0.792 0.468 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.576 0.756 ; 
        RECT 0.504 0.252 0.576 0.756 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
      LAYER M2 ; 
        RECT 0.292 0.54 0.652 0.612 ; 
      LAYER V1 ; 
        RECT 0.504 0.54 0.576 0.612 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
      LAYER M2 ; 
        RECT 0.072 0.396 0.328 0.468 ; 
      LAYER V1 ; 
        RECT 0.072 0.396 0.144 0.468 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.108 0.684 1.268 0.756 ; 
        RECT 1.152 0.396 1.224 0.756 ; 
      LAYER M2 ; 
        RECT 1.028 0.54 1.344 0.612 ; 
      LAYER V1 ; 
        RECT 1.152 0.54 1.224 0.612 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.36 0.54 1.588 0.612 ; 
        RECT 1.36 0.396 1.588 0.468 ; 
        RECT 1.36 0.396 1.432 0.612 ; 
      LAYER M2 ; 
        RECT 1.32 0.396 1.612 0.468 ; 
      LAYER V1 ; 
        RECT 1.44 0.396 1.512 0.468 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.252 1.084 0.324 ; 
        RECT 0.936 0.252 1.008 0.584 ; 
      LAYER M2 ; 
        RECT 0.848 0.252 1.112 0.324 ; 
      LAYER V1 ; 
        RECT 0.944 0.252 1.016 0.324 ; 
    END 
  END C 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.104 0.684 2.516 0.756 ; 
        RECT 2.444 0.108 2.516 0.756 ; 
        RECT 2.104 0.108 2.516 0.18 ; 
      LAYER M2 ; 
        RECT 1.836 0.396 2.516 0.468 ; 
      LAYER V1 ; 
        RECT 2.444 0.396 2.516 0.468 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.424 0.684 1.784 0.756 ; 
      RECT 1.712 0.252 1.784 0.756 ; 
      RECT 1.712 0.396 2.108 0.468 ; 
      RECT 1.26 0.252 1.784 0.324 ; 
      RECT 1.024 0.108 1.584 0.18 ; 
      RECT 0.792 0.684 0.952 0.756 ; 
      RECT 0.376 0.108 0.9 0.18 ; 
    LAYER M2 ; 
      RECT 0.828 0.684 1.764 0.756 ; 
    LAYER V1 ; 
      RECT 1.692 0.684 1.764 0.756 ; 
      RECT 0.828 0.684 0.9 0.756 ; 
  END 
END OA321x2_ASAP7_6t_SL 


MACRO OA322x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA322x1_ASAP7_6t_SL 0 0 ; 
  SIZE 2.592 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.148 0.252 2.236 0.548 ; 
        RECT 2.072 0.608 2.22 0.756 ; 
        RECT 2.148 0.252 2.22 0.756 ; 
        RECT 2.016 0.396 2.236 0.468 ; 
        RECT 2.088 0.252 2.236 0.468 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.608 2 0.756 ; 
        RECT 1.8 0.252 1.948 0.324 ; 
        RECT 1.8 0.252 1.872 0.756 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.436 0.252 1.7 0.324 ; 
        RECT 1.456 0.684 1.656 0.756 ; 
        RECT 1.584 0.252 1.656 0.756 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.832 0.54 1.068 0.612 ; 
        RECT 0.996 0.396 1.068 0.612 ; 
        RECT 0.836 0.396 1.068 0.468 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.14 0.396 1.444 0.468 ; 
        RECT 1.14 0.54 1.36 0.612 ; 
        RECT 1.14 0.396 1.212 0.612 ; 
    END 
  END B2 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.068 0.608 0.272 0.756 ; 
        RECT 0.068 0.252 0.216 0.756 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.488 0.396 0.712 0.468 ; 
        RECT 0.488 0.54 0.708 0.612 ; 
        RECT 0.488 0.396 0.56 0.612 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.592 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.32 0.684 2.524 0.756 ; 
        RECT 2.452 0.148 2.524 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 2.308 0.108 2.38 0.488 ; 
      RECT 2.104 0.108 2.38 0.18 ; 
      RECT 0.344 0.684 1.332 0.756 ; 
      RECT 0.344 0.404 0.416 0.756 ; 
      RECT 0.288 0.108 0.364 0.476 ; 
      RECT 0.128 0.108 0.364 0.18 ; 
      RECT 0.436 0.252 1.312 0.324 ; 
      RECT 0.436 0.16 0.508 0.324 ; 
      RECT 1.044 0.108 1.98 0.18 ; 
      RECT 0.772 0.108 0.92 0.18 ; 
    LAYER M2 ; 
      RECT 0.16 0.108 2.216 0.18 ; 
    LAYER V1 ; 
      RECT 2.124 0.108 2.196 0.18 ; 
      RECT 0.828 0.108 0.9 0.18 ; 
      RECT 0.18 0.108 0.252 0.18 ; 
  END 
END OA322x1_ASAP7_6t_SL 


MACRO OA322x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA322x2_ASAP7_6t_SL 0 0 ; 
  SIZE 2.808 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.1 0.108 2.248 0.26 ; 
        RECT 2.088 0.608 2.236 0.756 ; 
        RECT 2.164 0.108 2.236 0.756 ; 
        RECT 2.008 0.396 2.236 0.468 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.788 0.54 1.936 0.612 ; 
        RECT 1.788 0.252 1.936 0.324 ; 
        RECT 1.788 0.252 1.86 0.612 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.684 1.804 0.756 ; 
        RECT 1.584 0.252 1.656 0.756 ; 
        RECT 1.436 0.252 1.656 0.324 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.856 0.54 1.076 0.612 ; 
        RECT 1.004 0.396 1.076 0.612 ; 
        RECT 0.856 0.396 1.076 0.468 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.148 0.396 1.464 0.468 ; 
        RECT 1.148 0.54 1.444 0.612 ; 
        RECT 1.148 0.396 1.22 0.612 ; 
    END 
  END B2 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.064 0.608 0.272 0.756 ; 
        RECT 0.036 0.252 0.184 0.4 ; 
        RECT 0.064 0.252 0.136 0.756 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.488 0.396 0.712 0.468 ; 
        RECT 0.488 0.54 0.708 0.612 ; 
        RECT 0.488 0.396 0.56 0.612 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.808 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.808 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.316 0.608 2.464 0.756 ; 
        RECT 2.392 0.412 2.464 0.756 ; 
        RECT 2.316 0.312 2.392 0.484 ; 
        RECT 2.32 0.136 2.392 0.484 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 2.536 0.604 2.74 0.752 ; 
      RECT 2.668 0.108 2.74 0.752 ; 
      RECT 2.536 0.108 2.74 0.18 ; 
      RECT 0.344 0.684 1.368 0.756 ; 
      RECT 0.344 0.412 0.416 0.756 ; 
      RECT 0.292 0.108 0.364 0.484 ; 
      RECT 0.064 0.108 0.364 0.18 ; 
      RECT 0.436 0.252 1.312 0.324 ; 
      RECT 0.436 0.16 0.508 0.324 ; 
      RECT 1.044 0.108 2 0.18 ; 
      RECT 0.752 0.108 0.92 0.18 ; 
    LAYER M2 ; 
      RECT 0.14 0.108 2.732 0.18 ; 
    LAYER V1 ; 
      RECT 2.556 0.108 2.628 0.18 ; 
      RECT 0.828 0.108 0.9 0.18 ; 
      RECT 0.18 0.108 0.252 0.18 ; 
  END 
END OA322x2_ASAP7_6t_SL 


MACRO OA32x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA32x1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.856 0.548 1.004 0.696 ; 
        RECT 0.932 0.252 1.004 0.696 ; 
        RECT 0.856 0.252 1.004 0.4 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.636 0.548 0.784 0.696 ; 
        RECT 0.712 0.252 0.784 0.696 ; 
        RECT 0.636 0.252 0.784 0.4 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.492 0.252 0.564 0.604 ; 
        RECT 0.396 0.252 0.564 0.324 ; 
        RECT 0.34 0.108 0.488 0.256 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.36 1.224 0.696 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.516 0.528 1.664 0.608 ; 
        RECT 1.592 0.252 1.664 0.608 ; 
        RECT 1.44 0.252 1.664 0.4 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.092 0.108 0.24 0.18 ; 
        RECT 0.092 0.108 0.164 0.7 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.296 0.684 1.572 0.756 ; 
      RECT 1.296 0.224 1.368 0.756 ; 
      RECT 0.256 0.684 0.48 0.756 ; 
      RECT 0.256 0.396 0.328 0.756 ; 
      RECT 1.452 0.108 1.664 0.18 ; 
      RECT 0.612 0.108 1.148 0.18 ; 
    LAYER M2 ; 
      RECT 1.008 0.108 1.58 0.18 ; 
      RECT 0.376 0.684 1.576 0.756 ; 
    LAYER V1 ; 
      RECT 1.476 0.108 1.548 0.18 ; 
      RECT 1.476 0.684 1.548 0.756 ; 
      RECT 1.044 0.108 1.116 0.18 ; 
      RECT 0.396 0.684 0.468 0.756 ; 
  END 
END OA32x1_ASAP7_6t_SL 


MACRO OA32x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA32x2_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.072 0.548 1.22 0.696 ; 
        RECT 1.148 0.252 1.22 0.696 ; 
        RECT 1.072 0.252 1.22 0.4 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.852 0.548 1 0.696 ; 
        RECT 0.928 0.252 1 0.696 ; 
        RECT 0.852 0.252 1 0.4 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.708 0.252 0.78 0.676 ; 
        RECT 0.552 0.252 0.78 0.324 ; 
        RECT 0.552 0.108 0.696 0.324 ; 
        RECT 0.38 0.108 0.696 0.18 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.252 1.44 0.54 ; 
        RECT 1.292 0.252 1.44 0.4 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.76 0.528 1.908 0.756 ; 
        RECT 1.732 0.252 1.88 0.324 ; 
        RECT 1.732 0.252 1.804 0.608 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.54 0.448 0.612 ; 
        RECT 0.072 0.252 0.428 0.324 ; 
        RECT 0.072 0.54 0.22 0.756 ; 
        RECT 0.072 0.108 0.22 0.324 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.368 0.684 1.66 0.756 ; 
      RECT 1.512 0.224 1.584 0.756 ; 
      RECT 0.344 0.684 0.624 0.756 ; 
      RECT 0.548 0.396 0.62 0.756 ; 
      RECT 0.336 0.396 0.62 0.468 ; 
      RECT 1.668 0.108 1.88 0.18 ; 
      RECT 0.828 0.108 1.364 0.18 ; 
    LAYER M2 ; 
      RECT 1.24 0.108 1.784 0.18 ; 
      RECT 0.364 0.684 1.568 0.756 ; 
    LAYER V1 ; 
      RECT 1.692 0.108 1.764 0.18 ; 
      RECT 1.476 0.684 1.548 0.756 ; 
      RECT 1.26 0.108 1.332 0.18 ; 
      RECT 0.396 0.684 0.468 0.756 ; 
  END 
END OA32x2_ASAP7_6t_SL 


MACRO OA331x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA331x1_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.252 1.084 0.324 ; 
        RECT 0.896 0.684 1.044 0.756 ; 
        RECT 0.936 0.252 1.008 0.756 ; 
      LAYER M2 ; 
        RECT 0.82 0.252 1.204 0.324 ; 
      LAYER V1 ; 
        RECT 0.988 0.252 1.06 0.324 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.684 0.252 0.832 0.324 ; 
        RECT 0.648 0.684 0.796 0.756 ; 
        RECT 0.724 0.252 0.796 0.756 ; 
      LAYER M2 ; 
        RECT 0.524 0.396 0.988 0.468 ; 
      LAYER V1 ; 
        RECT 0.724 0.396 0.796 0.468 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.252 0.576 0.48 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
      LAYER M2 ; 
        RECT 0.304 0.252 0.692 0.324 ; 
      LAYER V1 ; 
        RECT 0.468 0.252 0.54 0.324 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.144 0.684 1.292 0.756 ; 
        RECT 1.144 0.396 1.216 0.756 ; 
      LAYER M2 ; 
        RECT 0.956 0.54 1.42 0.612 ; 
      LAYER V1 ; 
        RECT 1.144 0.54 1.216 0.612 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.336 0.396 1.484 0.468 ; 
        RECT 1.372 0.396 1.444 0.584 ; 
      LAYER M2 ; 
        RECT 1.172 0.396 1.648 0.468 ; 
      LAYER V1 ; 
        RECT 1.388 0.396 1.46 0.468 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.54 1.772 0.612 ; 
        RECT 1.584 0.424 1.656 0.612 ; 
      LAYER M2 ; 
        RECT 1.608 0.54 2.044 0.612 ; 
      LAYER V1 ; 
        RECT 1.692 0.54 1.764 0.612 ; 
    END 
  END B3 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.908 0.396 1.98 0.584 ; 
        RECT 1.808 0.396 1.98 0.468 ; 
      LAYER M2 ; 
        RECT 1.784 0.396 2.044 0.468 ; 
      LAYER V1 ; 
        RECT 1.876 0.396 1.948 0.468 ; 
    END 
  END C 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.684 0.252 0.756 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
      LAYER M2 ; 
        RECT 0.156 0.108 0.548 0.18 ; 
      LAYER V1 ; 
        RECT 0.18 0.108 0.252 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.456 0.684 2.124 0.756 ; 
      RECT 2.052 0.108 2.124 0.756 ; 
      RECT 1.808 0.108 2.124 0.18 ; 
      RECT 0.376 0.684 0.524 0.756 ; 
      RECT 0.376 0.54 0.448 0.756 ; 
      RECT 0.288 0.54 0.448 0.612 ; 
      RECT 0.288 0.376 0.36 0.612 ; 
      RECT 1.28 0.252 1.86 0.324 ; 
      RECT 0.576 0.108 1.572 0.18 ; 
    LAYER M2 ; 
      RECT 0.376 0.684 1.784 0.756 ; 
    LAYER V1 ; 
      RECT 1.692 0.684 1.764 0.756 ; 
      RECT 0.396 0.684 0.468 0.756 ; 
  END 
END OA331x1_ASAP7_6t_SL 


MACRO OA331x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA331x2_ASAP7_6t_SL 0 0 ; 
  SIZE 2.376 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.376 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.252 1.308 0.324 ; 
        RECT 1.152 0.252 1.224 0.652 ; 
      LAYER M2 ; 
        RECT 1.188 0.252 1.52 0.324 ; 
      LAYER V1 ; 
        RECT 1.188 0.252 1.26 0.324 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.9 0.252 1.048 0.324 ; 
        RECT 0.932 0.252 1.004 0.652 ; 
      LAYER M2 ; 
        RECT 0.836 0.54 1.116 0.612 ; 
      LAYER V1 ; 
        RECT 0.932 0.54 1.004 0.612 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.252 0.792 0.476 ; 
        RECT 0.644 0.252 0.792 0.324 ; 
      LAYER M2 ; 
        RECT 0.452 0.252 0.74 0.324 ; 
      LAYER V1 ; 
        RECT 0.668 0.252 0.74 0.324 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.344 0.396 1.456 0.468 ; 
        RECT 1.36 0.396 1.432 0.652 ; 
      LAYER M2 ; 
        RECT 1.36 0.396 1.648 0.468 ; 
      LAYER V1 ; 
        RECT 1.36 0.396 1.432 0.468 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.532 0.54 1.7 0.612 ; 
        RECT 1.588 0.424 1.66 0.612 ; 
      LAYER M2 ; 
        RECT 1.532 0.54 1.812 0.612 ; 
      LAYER V1 ; 
        RECT 1.552 0.54 1.624 0.612 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.54 2.136 0.612 ; 
        RECT 1.8 0.424 1.872 0.612 ; 
      LAYER M2 ; 
        RECT 1.936 0.54 2.22 0.612 ; 
      LAYER V1 ; 
        RECT 1.936 0.54 2.008 0.612 ; 
    END 
  END B3 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.996 0.396 2.168 0.468 ; 
      LAYER M2 ; 
        RECT 2 0.396 2.288 0.468 ; 
      LAYER V1 ; 
        RECT 2.076 0.396 2.148 0.468 ; 
    END 
  END C 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 0.488 0.18 ; 
        RECT 0.072 0.684 0.468 0.756 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
      LAYER M2 ; 
        RECT 0.072 0.108 1.024 0.18 ; 
      LAYER V1 ; 
        RECT 0.18 0.108 0.252 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.672 0.684 2.34 0.756 ; 
      RECT 2.268 0.108 2.34 0.756 ; 
      RECT 2.024 0.108 2.34 0.18 ; 
      RECT 0.592 0.684 0.74 0.756 ; 
      RECT 0.592 0.54 0.664 0.756 ; 
      RECT 0.504 0.54 0.664 0.612 ; 
      RECT 0.504 0.376 0.576 0.612 ; 
      RECT 1.496 0.252 2.076 0.324 ; 
      RECT 0.788 0.108 1.788 0.18 ; 
    LAYER M2 ; 
      RECT 0.612 0.684 1.864 0.756 ; 
    LAYER V1 ; 
      RECT 1.692 0.684 1.764 0.756 ; 
      RECT 0.612 0.684 0.684 0.756 ; 
  END 
END OA331x2_ASAP7_6t_SL 


MACRO OA332x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA332x1_ASAP7_6t_SL 0 0 ; 
  SIZE 3.024 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.636 0.404 0.8 0.476 ; 
        RECT 0.376 0.684 0.708 0.756 ; 
        RECT 0.636 0.232 0.708 0.756 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.272 0.54 0.564 0.612 ; 
        RECT 0.492 0.252 0.564 0.612 ; 
        RECT 0.376 0.252 0.564 0.324 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.684 0.22 0.756 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.684 0.996 0.756 ; 
        RECT 0.924 0.252 0.996 0.756 ; 
        RECT 0.848 0.252 0.996 0.324 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.068 0.684 1.352 0.756 ; 
        RECT 1.068 0.396 1.288 0.468 ; 
        RECT 1.068 0.396 1.14 0.756 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.24 0.54 1.648 0.612 ; 
        RECT 1.428 0.396 1.648 0.468 ; 
        RECT 1.428 0.396 1.5 0.612 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.368 0.54 2.528 0.612 ; 
        RECT 2.456 0.108 2.528 0.612 ; 
        RECT 2.32 0.108 2.528 0.18 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.78 0.54 2.12 0.612 ; 
        RECT 2.048 0.396 2.12 0.612 ; 
        RECT 1.78 0.396 2.12 0.468 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.024 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.024 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.804 0.684 2.952 0.756 ; 
        RECT 2.88 0.108 2.952 0.756 ; 
        RECT 2.752 0.108 2.952 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.476 0.684 2.672 0.756 ; 
      RECT 2.6 0.396 2.672 0.756 ; 
      RECT 2.196 0.252 2.268 0.756 ; 
      RECT 2.6 0.396 2.78 0.468 ; 
      RECT 1.928 0.252 2.268 0.324 ; 
      RECT 1.1 0.252 1.804 0.324 ; 
      RECT 1.732 0.108 1.804 0.324 ; 
      RECT 1.732 0.108 2.196 0.18 ; 
      RECT 0.772 0.108 1.568 0.18 ; 
      RECT 0.376 0.108 0.54 0.18 ; 
    LAYER M2 ; 
      RECT 0.396 0.108 0.936 0.18 ; 
    LAYER V1 ; 
      RECT 0.828 0.108 0.9 0.18 ; 
      RECT 0.396 0.108 0.468 0.18 ; 
  END 
END OA332x1_ASAP7_6t_SL 


MACRO OA332x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA332x2_ASAP7_6t_SL 0 0 ; 
  SIZE 3.24 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.636 0.404 0.8 0.476 ; 
        RECT 0.376 0.684 0.708 0.756 ; 
        RECT 0.636 0.232 0.708 0.756 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.272 0.54 0.564 0.612 ; 
        RECT 0.492 0.252 0.564 0.612 ; 
        RECT 0.376 0.252 0.564 0.324 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.684 0.22 0.756 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.684 0.996 0.756 ; 
        RECT 0.924 0.252 0.996 0.756 ; 
        RECT 0.828 0.252 0.996 0.324 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.068 0.684 1.352 0.756 ; 
        RECT 1.068 0.396 1.288 0.468 ; 
        RECT 1.068 0.396 1.14 0.756 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.24 0.54 1.648 0.612 ; 
        RECT 1.428 0.396 1.648 0.468 ; 
        RECT 1.428 0.396 1.5 0.612 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.368 0.54 2.528 0.612 ; 
        RECT 2.456 0.108 2.528 0.612 ; 
        RECT 2.32 0.108 2.528 0.18 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.78 0.54 2.12 0.612 ; 
        RECT 2.048 0.396 2.12 0.612 ; 
        RECT 1.78 0.396 2.12 0.468 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.24 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.24 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.804 0.684 3.168 0.756 ; 
        RECT 3.096 0.108 3.168 0.756 ; 
        RECT 2.808 0.108 3.168 0.18 ; 
        RECT 2.808 0.108 2.88 0.272 ; 
        RECT 2.804 0.592 2.876 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.476 0.684 2.7 0.756 ; 
      RECT 2.628 0.396 2.7 0.756 ; 
      RECT 2.196 0.252 2.268 0.756 ; 
      RECT 2.628 0.396 2.8 0.468 ; 
      RECT 1.928 0.252 2.268 0.324 ; 
      RECT 1.1 0.252 1.804 0.324 ; 
      RECT 1.732 0.108 1.804 0.324 ; 
      RECT 1.732 0.108 2.196 0.18 ; 
      RECT 0.772 0.108 1.568 0.18 ; 
      RECT 0.376 0.108 0.54 0.18 ; 
    LAYER M2 ; 
      RECT 0.396 0.108 0.936 0.18 ; 
    LAYER V1 ; 
      RECT 0.828 0.108 0.9 0.18 ; 
      RECT 0.396 0.108 0.468 0.18 ; 
  END 
END OA332x2_ASAP7_6t_SL 


MACRO OA333x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA333x1_ASAP7_6t_SL 0 0 ; 
  SIZE 3.456 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.736 0.54 2.884 0.612 ; 
        RECT 2.736 0.252 2.884 0.324 ; 
        RECT 2.736 0.252 2.808 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.516 0.252 2.664 0.612 ; 
        RECT 2.224 0.396 2.664 0.468 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.32 0.684 2.552 0.756 ; 
        RECT 2.32 0.54 2.392 0.756 ; 
        RECT 1.864 0.54 2.392 0.612 ; 
        RECT 1.864 0.396 2.084 0.468 ; 
        RECT 1.864 0.396 1.936 0.612 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.684 0.996 0.756 ; 
        RECT 0.924 0.252 0.996 0.756 ; 
        RECT 0.82 0.252 0.996 0.324 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.068 0.684 1.288 0.756 ; 
        RECT 1.068 0.396 1.288 0.468 ; 
        RECT 1.068 0.228 1.14 0.756 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.428 0.396 1.668 0.468 ; 
        RECT 1.24 0.54 1.648 0.612 ; 
        RECT 1.428 0.396 1.5 0.612 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.636 0.404 0.8 0.476 ; 
        RECT 0.376 0.684 0.708 0.756 ; 
        RECT 0.636 0.232 0.708 0.756 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.372 0.54 0.564 0.612 ; 
        RECT 0.492 0.252 0.564 0.612 ; 
        RECT 0.376 0.252 0.564 0.324 ; 
    END 
  END C2 
  PIN C3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END C3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.456 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.456 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 3.184 0.684 3.384 0.756 ; 
        RECT 3.312 0.108 3.384 0.756 ; 
        RECT 3.184 0.108 3.384 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 2.752 0.684 3.056 0.756 ; 
      RECT 2.984 0.528 3.056 0.756 ; 
      RECT 3.028 0.264 3.1 0.6 ; 
      RECT 2.984 0.108 3.056 0.336 ; 
      RECT 2.536 0.108 3.056 0.18 ; 
      RECT 1.252 0.252 2.412 0.324 ; 
      RECT 2.34 0.16 2.412 0.324 ; 
      RECT 1.252 0.16 1.324 0.324 ; 
      RECT 2.02 0.108 2.216 0.18 ; 
      RECT 1.456 0.684 2.196 0.756 ; 
      RECT 1.452 0.108 1.652 0.18 ; 
      RECT 0.772 0.108 0.956 0.18 ; 
      RECT 0.376 0.108 0.54 0.18 ; 
    LAYER M2 ; 
      RECT 2.084 0.108 2.72 0.18 ; 
      RECT 0.396 0.108 1.62 0.18 ; 
    LAYER V1 ; 
      RECT 2.556 0.108 2.628 0.18 ; 
      RECT 2.124 0.108 2.196 0.18 ; 
      RECT 1.476 0.108 1.548 0.18 ; 
      RECT 0.828 0.108 0.9 0.18 ; 
      RECT 0.396 0.108 0.468 0.18 ; 
  END 
END OA333x1_ASAP7_6t_SL 


MACRO OA333x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA333x2_ASAP7_6t_SL 0 0 ; 
  SIZE 3.672 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.736 0.54 2.884 0.612 ; 
        RECT 2.736 0.252 2.884 0.324 ; 
        RECT 2.736 0.252 2.808 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.516 0.252 2.664 0.612 ; 
        RECT 2.22 0.396 2.664 0.468 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.32 0.684 2.552 0.756 ; 
        RECT 2.32 0.54 2.392 0.756 ; 
        RECT 1.864 0.54 2.392 0.612 ; 
        RECT 1.864 0.396 2.088 0.468 ; 
        RECT 1.864 0.396 1.936 0.612 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.684 0.996 0.756 ; 
        RECT 0.924 0.252 0.996 0.756 ; 
        RECT 0.82 0.252 0.996 0.324 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.068 0.684 1.288 0.756 ; 
        RECT 1.068 0.396 1.288 0.468 ; 
        RECT 1.068 0.228 1.14 0.756 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.24 0.54 1.648 0.612 ; 
        RECT 1.428 0.396 1.648 0.468 ; 
        RECT 1.428 0.396 1.5 0.612 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.636 0.404 0.8 0.476 ; 
        RECT 0.376 0.684 0.708 0.756 ; 
        RECT 0.636 0.232 0.708 0.756 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.364 0.54 0.564 0.612 ; 
        RECT 0.492 0.252 0.564 0.612 ; 
        RECT 0.376 0.252 0.564 0.324 ; 
    END 
  END C2 
  PIN C3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.684 0.252 0.756 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END C3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 3.672 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.672 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 3.184 0.684 3.384 0.756 ; 
        RECT 3.312 0.108 3.384 0.756 ; 
        RECT 3.184 0.108 3.384 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 2.752 0.684 3.08 0.756 ; 
      RECT 3.008 0.528 3.08 0.756 ; 
      RECT 3.028 0.256 3.1 0.6 ; 
      RECT 3.008 0.108 3.08 0.328 ; 
      RECT 2.536 0.108 3.08 0.18 ; 
      RECT 1.252 0.252 2.412 0.324 ; 
      RECT 2.34 0.16 2.412 0.324 ; 
      RECT 1.252 0.16 1.324 0.324 ; 
      RECT 2.02 0.108 2.216 0.18 ; 
      RECT 1.456 0.684 2.196 0.756 ; 
      RECT 1.452 0.108 1.652 0.18 ; 
      RECT 0.772 0.108 0.956 0.18 ; 
      RECT 0.376 0.108 0.54 0.18 ; 
    LAYER M2 ; 
      RECT 2.084 0.108 2.72 0.18 ; 
      RECT 0.396 0.108 1.62 0.18 ; 
    LAYER V1 ; 
      RECT 2.556 0.108 2.628 0.18 ; 
      RECT 2.124 0.108 2.196 0.18 ; 
      RECT 1.476 0.108 1.548 0.18 ; 
      RECT 0.828 0.108 0.9 0.18 ; 
      RECT 0.396 0.108 0.468 0.18 ; 
  END 
END OA333x2_ASAP7_6t_SL 


MACRO OA33x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA33x1_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.608 1.008 0.756 ; 
        RECT 0.936 0.252 1.008 0.756 ; 
        RECT 0.748 0.252 1.008 0.324 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.108 0.252 1.268 0.324 ; 
        RECT 1.108 0.54 1.26 0.612 ; 
        RECT 1.152 0.252 1.224 0.612 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.548 0.396 0.812 0.468 ; 
        RECT 0.548 0.684 0.704 0.756 ; 
        RECT 0.548 0.184 0.62 0.756 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.12 0.684 1.432 0.756 ; 
        RECT 1.36 0.424 1.432 0.756 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.504 0.684 1.832 0.756 ; 
        RECT 1.504 0.396 1.668 0.468 ; 
        RECT 1.504 0.396 1.576 0.756 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.94 0.684 2.096 0.756 ; 
        RECT 1.94 0.396 2.088 0.468 ; 
        RECT 1.94 0.396 2.012 0.756 ; 
    END 
  END B3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.284 0.572 0.448 0.644 ; 
        RECT 0.284 0.252 0.448 0.324 ; 
        RECT 0.08 0.684 0.356 0.756 ; 
        RECT 0.284 0.252 0.356 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.704 0.54 1.868 0.612 ; 
      RECT 1.796 0.252 1.868 0.612 ; 
      RECT 1.412 0.252 2.016 0.324 ; 
      RECT 1.888 0.108 2.016 0.324 ; 
      RECT 1.888 0.108 2.088 0.18 ; 
      RECT 0.072 0.108 0.144 0.496 ; 
      RECT 0.072 0.108 0.292 0.18 ; 
      RECT 0.804 0.108 1.764 0.18 ; 
    LAYER M2 ; 
      RECT 0.1 0.108 2.052 0.18 ; 
    LAYER V1 ; 
      RECT 1.908 0.108 1.98 0.18 ; 
      RECT 0.18 0.108 0.252 0.18 ; 
  END 
END OA33x1_ASAP7_6t_SL 


MACRO OA33x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA33x2_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.608 1.008 0.756 ; 
        RECT 0.936 0.252 1.008 0.756 ; 
        RECT 0.748 0.252 1.008 0.324 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.108 0.252 1.268 0.324 ; 
        RECT 1.108 0.54 1.26 0.612 ; 
        RECT 1.152 0.252 1.224 0.612 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.548 0.396 0.792 0.468 ; 
        RECT 0.548 0.608 0.704 0.756 ; 
        RECT 0.548 0.212 0.62 0.756 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.12 0.684 1.432 0.756 ; 
        RECT 1.36 0.424 1.432 0.756 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.504 0.684 1.782 0.756 ; 
        RECT 1.504 0.396 1.668 0.468 ; 
        RECT 1.504 0.396 1.576 0.756 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.952 0.54 2.124 0.756 ; 
        RECT 2.024 0.396 2.096 0.756 ; 
    END 
  END B3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.284 0.572 0.448 0.644 ; 
        RECT 0.356 0.232 0.428 0.448 ; 
        RECT 0.08 0.684 0.356 0.756 ; 
        RECT 0.284 0.376 0.356 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.704 0.54 1.868 0.612 ; 
      RECT 1.796 0.252 1.868 0.612 ; 
      RECT 1.412 0.252 1.988 0.324 ; 
      RECT 1.896 0.108 1.988 0.324 ; 
      RECT 1.896 0.108 2.088 0.18 ; 
      RECT 0.072 0.108 0.144 0.496 ; 
      RECT 0.072 0.108 0.272 0.184 ; 
      RECT 0.804 0.108 1.764 0.18 ; 
    LAYER M2 ; 
      RECT 0.1 0.108 2.052 0.18 ; 
    LAYER V1 ; 
      RECT 1.908 0.108 1.98 0.18 ; 
      RECT 0.18 0.108 0.252 0.18 ; 
  END 
END OA33x2_ASAP7_6t_SL 


MACRO OAI211xp33_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI211xp33_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.388 0.576 0.584 ; 
      LAYER M2 ; 
        RECT 0.384 0.396 0.68 0.468 ; 
      LAYER V1 ; 
        RECT 0.504 0.396 0.576 0.468 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.064 0.684 0.216 0.756 ; 
        RECT 0.144 0.252 0.216 0.756 ; 
        RECT 0.064 0.252 0.216 0.324 ; 
      LAYER M2 ; 
        RECT 0.072 0.54 0.46 0.612 ; 
      LAYER V1 ; 
        RECT 0.144 0.54 0.216 0.612 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.54 0.92 0.612 ; 
        RECT 0.72 0.252 0.792 0.612 ; 
        RECT 0.628 0.252 0.792 0.324 ; 
      LAYER M2 ; 
        RECT 0.54 0.252 0.892 0.324 ; 
      LAYER V1 ; 
        RECT 0.652 0.252 0.724 0.324 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.044 0.304 1.116 0.568 ; 
        RECT 0.936 0.304 1.116 0.376 ; 
        RECT 0.936 0.108 1.008 0.376 ; 
        RECT 0.828 0.108 1.008 0.18 ; 
      LAYER M2 ; 
        RECT 0.872 0.396 1.18 0.468 ; 
      LAYER V1 ; 
        RECT 1.044 0.396 1.116 0.468 ; 
    END 
  END C 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.684 1.26 0.756 ; 
        RECT 1.188 0.108 1.26 0.756 ; 
        RECT 1.112 0.108 1.26 0.18 ; 
        RECT 0.288 0.252 0.452 0.324 ; 
        RECT 0.288 0.252 0.36 0.756 ; 
      LAYER M2 ; 
        RECT 0.624 0.684 1.232 0.756 ; 
      LAYER V1 ; 
        RECT 1.044 0.684 1.116 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.108 0.704 0.18 ; 
  END 
END OAI211xp33_ASAP7_6t_SL 


MACRO OAI211xp67b_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI211xp67b_ASAP7_6t_SL 0 0 ; 
  SIZE 2.592 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.592 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.636 0.396 0.952 0.468 ; 
        RECT 0.636 0.684 0.936 0.756 ; 
        RECT 0.636 0.252 0.936 0.324 ; 
        RECT 0.636 0.252 0.708 0.756 ; 
      LAYER M2 ; 
        RECT 0.672 0.396 0.928 0.468 ; 
      LAYER V1 ; 
        RECT 0.808 0.396 0.88 0.468 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.492 0.468 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
      LAYER M2 ; 
        RECT 0.072 0.252 0.444 0.324 ; 
      LAYER V1 ; 
        RECT 0.072 0.252 0.144 0.324 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.256 0.684 1.476 0.756 ; 
        RECT 1.256 0.396 1.476 0.468 ; 
        RECT 1.256 0.396 1.328 0.756 ; 
      LAYER M2 ; 
        RECT 1.16 0.54 1.416 0.612 ; 
      LAYER V1 ; 
        RECT 1.256 0.54 1.328 0.612 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.104 0.684 2.256 0.756 ; 
        RECT 2.184 0.396 2.256 0.756 ; 
        RECT 2.076 0.396 2.256 0.468 ; 
      LAYER M2 ; 
        RECT 2.076 0.54 2.336 0.612 ; 
      LAYER V1 ; 
        RECT 2.184 0.54 2.256 0.612 ; 
    END 
  END C 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.332 0.684 2.524 0.756 ; 
        RECT 2.332 0.252 2.412 0.756 ; 
        RECT 2.076 0.252 2.412 0.324 ; 
        RECT 1.672 0.684 1.98 0.756 ; 
        RECT 0.376 0.684 0.524 0.756 ; 
      LAYER M2 ; 
        RECT 0.396 0.684 2.48 0.756 ; 
      LAYER V1 ; 
        RECT 0.396 0.684 0.468 0.756 ; 
        RECT 1.692 0.684 1.764 0.756 ; 
        RECT 2.34 0.684 2.412 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.152 0.252 1.796 0.324 ; 
      RECT 1.152 0.108 1.224 0.324 ; 
      RECT 0.376 0.108 1.224 0.18 ; 
      RECT 1.444 0.108 2.432 0.18 ; 
  END 
END OAI211xp67b_ASAP7_6t_SL 


MACRO OAI21xp25_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21xp25_ASAP7_6t_SL 0 0 ; 
  SIZE 1.08 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.344 0.4 0.596 0.472 ; 
        RECT 0.344 0.252 0.576 0.324 ; 
        RECT 0.344 0.608 0.492 0.756 ; 
        RECT 0.344 0.252 0.416 0.756 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.252 0.22 0.324 ; 
        RECT 0.072 0.252 0.144 0.756 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.54 0.868 0.612 ; 
        RECT 0.72 0.252 0.868 0.324 ; 
        RECT 0.72 0.252 0.792 0.612 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.08 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.08 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.684 1.044 0.756 ; 
        RECT 0.972 0.108 1.044 0.756 ; 
        RECT 0.808 0.108 1.044 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.108 0.684 0.18 ; 
  END 
END OAI21xp25_ASAP7_6t_SL 


MACRO OAI21xp5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21xp5_ASAP7_6t_SL 0 0 ; 
  SIZE 1.08 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.344 0.4 0.576 0.472 ; 
        RECT 0.344 0.252 0.576 0.324 ; 
        RECT 0.344 0.4 0.492 0.756 ; 
        RECT 0.344 0.252 0.416 0.756 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.592 0.272 0.756 ; 
        RECT 0.072 0.252 0.244 0.324 ; 
        RECT 0.072 0.252 0.144 0.756 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.54 0.868 0.612 ; 
        RECT 0.72 0.252 0.868 0.324 ; 
        RECT 0.72 0.252 0.792 0.612 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.08 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.08 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.684 1.044 0.756 ; 
        RECT 0.972 0.108 1.044 0.756 ; 
        RECT 0.808 0.108 1.044 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.108 0.684 0.18 ; 
  END 
END OAI21xp5_ASAP7_6t_SL 


MACRO OAI21xp5b_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21xp5b_ASAP7_6t_SL 0 0 ; 
  SIZE 1.08 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.064 0.684 0.212 0.756 ; 
        RECT 0.14 0.252 0.212 0.756 ; 
        RECT 0.064 0.252 0.212 0.324 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.58 0.252 0.784 0.612 ; 
        RECT 0.488 0.4 0.784 0.472 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.856 0.684 1.004 0.756 ; 
        RECT 0.856 0.108 1.004 0.18 ; 
        RECT 0.856 0.108 0.928 0.756 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.08 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.08 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.284 0.684 0.708 0.756 ; 
        RECT 0.284 0.252 0.456 0.324 ; 
        RECT 0.284 0.252 0.356 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.108 0.704 0.18 ; 
  END 
END OAI21xp5b_ASAP7_6t_SL 


MACRO OAI221xp33_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI221xp33_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.056 0.252 1.204 0.324 ; 
        RECT 1.016 0.396 1.128 0.728 ; 
        RECT 1.056 0.252 1.128 0.728 ; 
        RECT 0.936 0.396 1.128 0.468 ; 
      LAYER M2 ; 
        RECT 0.884 0.252 1.312 0.324 ; 
      LAYER V1 ; 
        RECT 1.1 0.252 1.172 0.324 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.328 0.252 1.476 0.4 ; 
        RECT 1.228 0.684 1.448 0.756 ; 
        RECT 1.376 0.252 1.448 0.756 ; 
        RECT 1.228 0.54 1.448 0.612 ; 
      LAYER M2 ; 
        RECT 0.944 0.684 1.36 0.756 ; 
      LAYER V1 ; 
        RECT 1.26 0.684 1.332 0.756 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.036 0.608 0.188 0.756 ; 
        RECT 0.064 0.536 0.188 0.756 ; 
        RECT 0.036 0.252 0.188 0.4 ; 
        RECT 0.064 0.252 0.136 0.756 ; 
      LAYER M2 ; 
        RECT 0.068 0.54 0.512 0.612 ; 
      LAYER V1 ; 
        RECT 0.088 0.54 0.16 0.612 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.404 0.396 0.588 0.468 ; 
        RECT 0.404 0.396 0.48 0.584 ; 
      LAYER M2 ; 
        RECT 0.18 0.396 0.608 0.468 ; 
      LAYER V1 ; 
        RECT 0.496 0.396 0.568 0.468 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.54 0.868 0.612 ; 
        RECT 0.636 0.252 0.868 0.324 ; 
        RECT 0.72 0.252 0.792 0.612 ; 
      LAYER M2 ; 
        RECT 0.676 0.54 1.092 0.612 ; 
      LAYER V1 ; 
        RECT 0.728 0.54 0.8 0.612 ; 
    END 
  END C 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.26 0.684 0.9 0.756 ; 
        RECT 0.26 0.252 0.48 0.324 ; 
        RECT 0.26 0.252 0.332 0.756 ; 
      LAYER M2 ; 
        RECT 0.228 0.684 0.804 0.756 ; 
      LAYER V1 ; 
        RECT 0.396 0.684 0.468 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.828 0.108 1.448 0.18 ; 
      RECT 0.16 0.108 0.684 0.18 ; 
  END 
END OAI221xp33_ASAP7_6t_SL 


MACRO OAI221xp33f_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI221xp33f_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.684 1.172 0.756 ; 
        RECT 1.1 0.252 1.172 0.756 ; 
        RECT 0.936 0.396 1.172 0.468 ; 
        RECT 0.952 0.252 1.172 0.324 ; 
      LAYER M2 ; 
        RECT 0.94 0.252 1.216 0.324 ; 
      LAYER V1 ; 
        RECT 1.016 0.252 1.088 0.324 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.292 0.68 1.44 0.752 ; 
        RECT 1.368 0.252 1.44 0.752 ; 
        RECT 1.292 0.252 1.44 0.324 ; 
      LAYER M2 ; 
        RECT 1.164 0.396 1.44 0.468 ; 
      LAYER V1 ; 
        RECT 1.368 0.396 1.44 0.468 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.064 0.536 0.212 0.756 ; 
        RECT 0.064 0.28 0.136 0.756 ; 
      LAYER M2 ; 
        RECT 0.064 0.396 0.34 0.468 ; 
      LAYER V1 ; 
        RECT 0.064 0.396 0.136 0.468 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.456 0.54 0.604 0.612 ; 
        RECT 0.504 0.424 0.576 0.612 ; 
      LAYER M2 ; 
        RECT 0.44 0.54 0.696 0.612 ; 
      LAYER V1 ; 
        RECT 0.484 0.54 0.556 0.612 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.536 0.872 0.612 ; 
        RECT 0.72 0.252 0.792 0.612 ; 
        RECT 0.64 0.252 0.792 0.324 ; 
      LAYER M2 ; 
        RECT 0.628 0.396 0.904 0.468 ; 
      LAYER V1 ; 
        RECT 0.72 0.396 0.792 0.468 ; 
    END 
  END C 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.284 0.684 0.9 0.756 ; 
        RECT 0.284 0.252 0.468 0.324 ; 
        RECT 0.284 0.252 0.356 0.756 ; 
      LAYER M2 ; 
        RECT 0.284 0.252 0.776 0.324 ; 
      LAYER V1 ; 
        RECT 0.356 0.252 0.428 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.828 0.108 1.332 0.18 ; 
      RECT 0.16 0.108 0.684 0.18 ; 
  END 
END OAI221xp33f_ASAP7_6t_SL 


MACRO OAI222xp33_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI222xp33_ASAP7_6t_SL 0 0 ; 
  SIZE 2.16 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.16 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.036 0.528 0.184 0.756 ; 
        RECT 0.072 0.28 0.144 0.756 ; 
      LAYER M2 ; 
        RECT 0.072 0.396 0.352 0.468 ; 
      LAYER V1 ; 
        RECT 0.072 0.396 0.144 0.468 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.512 0.396 0.628 0.468 ; 
        RECT 0.436 0.54 0.584 0.612 ; 
        RECT 0.512 0.396 0.584 0.612 ; 
      LAYER M2 ; 
        RECT 0.412 0.54 0.748 0.612 ; 
      LAYER V1 ; 
        RECT 0.46 0.54 0.532 0.612 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.2 0.54 1.42 0.612 ; 
        RECT 1.348 0.396 1.42 0.612 ; 
        RECT 1.136 0.396 1.42 0.468 ; 
      LAYER M2 ; 
        RECT 1.148 0.54 1.484 0.612 ; 
      LAYER V1 ; 
        RECT 1.252 0.54 1.324 0.612 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.728 0.54 0.948 0.612 ; 
        RECT 0.728 0.396 0.948 0.468 ; 
        RECT 0.728 0.396 0.8 0.612 ; 
      LAYER M2 ; 
        RECT 0.656 0.396 1.04 0.468 ; 
      LAYER V1 ; 
        RECT 0.8 0.396 0.872 0.468 ; 
    END 
  END B2 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.656 0.608 1.804 0.756 ; 
        RECT 1.732 0.252 1.804 0.756 ; 
        RECT 1.564 0.396 1.804 0.468 ; 
        RECT 1.584 0.252 1.804 0.324 ; 
      LAYER M2 ; 
        RECT 1.46 0.396 1.844 0.468 ; 
      LAYER V1 ; 
        RECT 1.684 0.396 1.756 0.468 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.876 0.608 2.096 0.756 ; 
        RECT 2.024 0.108 2.096 0.756 ; 
        RECT 1.884 0.108 2.096 0.256 ; 
      LAYER M2 ; 
        RECT 1.62 0.252 2.096 0.324 ; 
      LAYER V1 ; 
        RECT 2.024 0.252 2.096 0.324 ; 
    END 
  END C2 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.256 0.684 1.352 0.756 ; 
        RECT 0.256 0.252 0.468 0.324 ; 
        RECT 0.256 0.252 0.328 0.756 ; 
      LAYER M2 ; 
        RECT 0.276 0.252 0.748 0.324 ; 
      LAYER V1 ; 
        RECT 0.324 0.252 0.396 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.796 0.252 1.44 0.324 ; 
      RECT 1.368 0.108 1.44 0.324 ; 
      RECT 1.368 0.108 1.784 0.18 ; 
      RECT 0.16 0.108 1.136 0.18 ; 
  END 
END OAI222xp33_ASAP7_6t_SL 


MACRO OAI22xp5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI22xp5_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.124 0.608 0.272 0.756 ; 
        RECT 0.124 0.252 0.272 0.4 ; 
        RECT 0.124 0.252 0.196 0.756 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.42 0.4 0.572 0.472 ; 
        RECT 0.344 0.608 0.492 0.756 ; 
        RECT 0.42 0.252 0.492 0.756 ; 
        RECT 0.344 0.252 0.492 0.4 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.684 1.176 0.756 ; 
        RECT 1.104 0.252 1.176 0.756 ; 
        RECT 1.024 0.252 1.176 0.4 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.58 0.608 0.78 0.756 ; 
        RECT 0.708 0.252 0.78 0.756 ; 
        RECT 0.608 0.252 0.78 0.324 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.852 0.232 0.924 0.644 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.992 0.108 1.14 0.18 ; 
      RECT 0.16 0.108 0.704 0.18 ; 
    LAYER M2 ; 
      RECT 0.592 0.108 1.136 0.18 ; 
    LAYER V1 ; 
      RECT 1.044 0.108 1.116 0.18 ; 
      RECT 0.612 0.108 0.684 0.18 ; 
  END 
END OAI22xp5_ASAP7_6t_SL 


MACRO OAI311xp33_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI311xp33_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.54 0.868 0.612 ; 
        RECT 0.72 0.376 0.792 0.612 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.576 0.756 ; 
        RECT 0.504 0.252 0.576 0.756 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.404 0.372 0.476 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A3 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.252 1.008 0.488 ; 
        RECT 0.86 0.252 1.008 0.324 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.148 0.54 1.296 0.612 ; 
        RECT 1.224 0.252 1.296 0.612 ; 
        RECT 1.14 0.252 1.296 0.324 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.792 0.684 1.44 0.756 ; 
        RECT 1.368 0.108 1.44 0.756 ; 
        RECT 1.22 0.108 1.44 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.108 0.92 0.18 ; 
  END 
END OAI311xp33_ASAP7_6t_SL 


MACRO OAI31x1f_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI31x1f_ASAP7_6t_SL 0 0 ; 
  SIZE 2.808 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.536 0.54 2.756 0.612 ; 
        RECT 2.684 0.396 2.756 0.612 ; 
        RECT 1.92 0.396 2.756 0.468 ; 
        RECT 2.32 0.108 2.468 0.18 ; 
        RECT 2.32 0.108 2.392 0.468 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.092 0.396 1.796 0.468 ; 
        RECT 1.092 0.684 1.312 0.756 ; 
        RECT 1.092 0.252 1.312 0.324 ; 
        RECT 1.092 0.252 1.164 0.756 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.372 0.468 ; 
        RECT 0.072 0.252 0.292 0.324 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.252 0.144 0.756 ; 
    END 
  END A3 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.616 0.396 0.788 0.468 ; 
        RECT 0.468 0.54 0.688 0.612 ; 
        RECT 0.616 0.252 0.688 0.612 ; 
        RECT 0.484 0.252 0.688 0.324 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.808 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.808 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.828 0.252 2.652 0.324 ; 
      LAYER M1 ; 
        RECT 2.516 0.252 2.696 0.324 ; 
        RECT 0.804 0.684 1.02 0.756 ; 
        RECT 0.948 0.252 1.02 0.756 ; 
        RECT 0.828 0.252 1.02 0.324 ; 
      LAYER V1 ; 
        RECT 0.928 0.252 1 0.324 ; 
        RECT 2.56 0.252 2.632 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 2.104 0.684 2.652 0.756 ; 
      RECT 1.456 0.54 2.412 0.612 ; 
      RECT 0.16 0.108 2.216 0.18 ; 
      RECT 1.632 0.684 1.788 0.756 ; 
      RECT 0.372 0.684 0.52 0.756 ; 
    LAYER M2 ; 
      RECT 0.376 0.684 1.788 0.756 ; 
    LAYER V1 ; 
      RECT 1.692 0.684 1.764 0.756 ; 
      RECT 0.396 0.684 0.468 0.756 ; 
  END 
END OAI31x1f_ASAP7_6t_SL 


MACRO OAI31xp5f_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI31xp5f_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.616 0.54 0.78 0.612 ; 
        RECT 0.708 0.252 0.78 0.612 ; 
        RECT 0.616 0.252 0.78 0.324 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.42 0.4 0.564 0.472 ; 
        RECT 0.344 0.608 0.492 0.756 ; 
        RECT 0.42 0.252 0.492 0.756 ; 
        RECT 0.344 0.252 0.492 0.324 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.248 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A3 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.88 0.54 1.028 0.612 ; 
        RECT 0.956 0.252 1.028 0.612 ; 
        RECT 0.88 0.252 1.028 0.324 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.732 0.684 1.224 0.756 ; 
        RECT 1.152 0.224 1.224 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.372 0.108 0.956 0.18 ; 
  END 
END OAI31xp5f_ASAP7_6t_SL 


MACRO OAI321xp33_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI321xp33_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.648 0.252 0.796 0.4 ; 
        RECT 0.72 0.252 0.792 0.584 ; 
      LAYER M2 ; 
        RECT 0.632 0.396 0.888 0.468 ; 
      LAYER V1 ; 
        RECT 0.72 0.396 0.792 0.468 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.576 0.756 ; 
        RECT 0.504 0.252 0.576 0.756 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
      LAYER M2 ; 
        RECT 0.388 0.54 0.652 0.612 ; 
      LAYER V1 ; 
        RECT 0.504 0.54 0.576 0.612 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
      LAYER M2 ; 
        RECT 0.072 0.252 0.42 0.324 ; 
      LAYER V1 ; 
        RECT 0.072 0.252 0.144 0.324 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.396 1.3 0.468 ; 
        RECT 1.108 0.684 1.268 0.756 ; 
        RECT 1.152 0.396 1.224 0.756 ; 
      LAYER M2 ; 
        RECT 1.072 0.396 1.388 0.468 ; 
      LAYER V1 ; 
        RECT 1.172 0.396 1.244 0.468 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.336 0.54 1.512 0.612 ; 
        RECT 1.44 0.424 1.512 0.612 ; 
      LAYER M2 ; 
        RECT 1.344 0.54 1.612 0.612 ; 
      LAYER V1 ; 
        RECT 1.344 0.54 1.416 0.612 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.252 1.084 0.324 ; 
        RECT 0.936 0.252 1.008 0.584 ; 
      LAYER M2 ; 
        RECT 0.848 0.252 1.112 0.324 ; 
      LAYER V1 ; 
        RECT 0.944 0.252 1.016 0.324 ; 
    END 
  END C 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.424 0.684 1.656 0.756 ; 
        RECT 1.584 0.252 1.656 0.756 ; 
        RECT 1.26 0.252 1.656 0.324 ; 
        RECT 0.792 0.684 0.952 0.756 ; 
      LAYER M2 ; 
        RECT 0.828 0.684 1.548 0.756 ; 
      LAYER V1 ; 
        RECT 0.828 0.684 0.9 0.756 ; 
        RECT 1.476 0.684 1.548 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.044 0.108 1.584 0.18 ; 
      RECT 0.396 0.108 0.9 0.18 ; 
  END 
END OAI321xp33_ASAP7_6t_SL 


MACRO OAI322xp33_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI322xp33_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.636 0.396 0.784 0.468 ; 
        RECT 0.636 0.396 0.708 0.62 ; 
      LAYER M2 ; 
        RECT 0.564 0.396 0.88 0.468 ; 
      LAYER V1 ; 
        RECT 0.68 0.396 0.752 0.468 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.82 0.54 1.008 0.612 ; 
        RECT 0.936 0.424 1.008 0.612 ; 
      LAYER M2 ; 
        RECT 0.808 0.54 1.08 0.612 ; 
      LAYER V1 ; 
        RECT 0.828 0.54 0.9 0.612 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.184 0.252 1.332 0.324 ; 
        RECT 1.12 0.684 1.268 0.756 ; 
        RECT 1.184 0.252 1.256 0.508 ; 
        RECT 1.152 0.44 1.224 0.756 ; 
      LAYER M2 ; 
        RECT 1.084 0.252 1.448 0.324 ; 
      LAYER V1 ; 
        RECT 1.208 0.252 1.28 0.324 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.564 0.756 ; 
        RECT 0.492 0.396 0.564 0.756 ; 
        RECT 0.336 0.396 0.564 0.468 ; 
      LAYER M2 ; 
        RECT 0.304 0.54 0.612 0.612 ; 
      LAYER V1 ; 
        RECT 0.492 0.54 0.564 0.612 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.252 0.284 0.324 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.252 0.144 0.756 ; 
      LAYER M2 ; 
        RECT 0.072 0.252 0.388 0.324 ; 
      LAYER V1 ; 
        RECT 0.146 0.252 0.218 0.324 ; 
    END 
  END B2 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.552 0.54 1.72 0.612 ; 
        RECT 1.648 0.424 1.72 0.612 ; 
      LAYER M2 ; 
        RECT 1.512 0.54 1.792 0.612 ; 
      LAYER V1 ; 
        RECT 1.56 0.54 1.632 0.612 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.684 1.516 0.756 ; 
        RECT 1.368 0.396 1.516 0.468 ; 
        RECT 1.368 0.396 1.44 0.756 ; 
      LAYER M2 ; 
        RECT 1.304 0.396 1.6 0.468 ; 
      LAYER V1 ; 
        RECT 1.404 0.396 1.476 0.468 ; 
    END 
  END C2 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.652 0.684 1.872 0.756 ; 
        RECT 1.8 0.252 1.872 0.756 ; 
        RECT 1.476 0.252 1.872 0.324 ; 
        RECT 0.776 0.684 0.996 0.756 ; 
      LAYER M2 ; 
        RECT 0.808 0.684 1.784 0.756 ; 
      LAYER V1 ; 
        RECT 0.828 0.684 0.9 0.756 ; 
        RECT 1.692 0.684 1.764 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.408 0.252 1.068 0.324 ; 
      RECT 0.408 0.108 0.48 0.324 ; 
      RECT 0.18 0.108 0.684 0.18 ; 
      RECT 0.828 0.108 1.8 0.18 ; 
  END 
END OAI322xp33_ASAP7_6t_SL 


MACRO OAI322xp33b_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI322xp33b_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.648 0.396 0.812 0.468 ; 
        RECT 0.648 0.396 0.72 0.636 ; 
      LAYER M2 ; 
        RECT 0.6 0.396 0.856 0.468 ; 
      LAYER V1 ; 
        RECT 0.68 0.396 0.752 0.468 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.888 0.54 1.044 0.612 ; 
        RECT 0.936 0.424 1.008 0.612 ; 
      LAYER M2 ; 
        RECT 0.828 0.54 1.132 0.612 ; 
      LAYER V1 ; 
        RECT 0.964 0.54 1.036 0.612 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.384 1.224 0.728 ; 
      LAYER M2 ; 
        RECT 0.988 0.396 1.244 0.468 ; 
      LAYER V1 ; 
        RECT 1.152 0.396 1.224 0.468 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.576 0.756 ; 
        RECT 0.504 0.396 0.576 0.756 ; 
        RECT 0.264 0.396 0.576 0.472 ; 
      LAYER M2 ; 
        RECT 0.356 0.54 0.684 0.612 ; 
      LAYER V1 ; 
        RECT 0.504 0.54 0.576 0.612 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.252 0.292 0.324 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.252 0.144 0.756 ; 
      LAYER M2 ; 
        RECT 0.072 0.252 0.36 0.324 ; 
      LAYER V1 ; 
        RECT 0.16 0.252 0.232 0.324 ; 
    END 
  END B2 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.732 0.68 1.88 0.756 ; 
        RECT 1.732 0.396 1.88 0.468 ; 
        RECT 1.732 0.28 1.804 0.756 ; 
      LAYER M2 ; 
        RECT 1.616 0.54 1.872 0.612 ; 
      LAYER V1 ; 
        RECT 1.732 0.54 1.804 0.612 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.336 0.396 1.484 0.468 ; 
        RECT 1.376 0.396 1.448 0.568 ; 
      LAYER M2 ; 
        RECT 1.368 0.396 1.624 0.468 ; 
      LAYER V1 ; 
        RECT 1.392 0.396 1.464 0.468 ; 
    END 
  END C2 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.412 0.684 1.656 0.756 ; 
        RECT 1.584 0.252 1.656 0.756 ; 
        RECT 1.436 0.252 1.656 0.324 ; 
        RECT 0.808 0.684 1.024 0.756 ; 
      LAYER M2 ; 
        RECT 0.828 0.684 1.548 0.756 ; 
      LAYER V1 ; 
        RECT 0.828 0.684 0.9 0.756 ; 
        RECT 1.476 0.684 1.548 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.416 0.252 1.096 0.324 ; 
      RECT 0.416 0.108 0.488 0.324 ; 
      RECT 0.18 0.108 0.684 0.18 ; 
      RECT 0.828 0.108 1.784 0.18 ; 
  END 
END OAI322xp33b_ASAP7_6t_SL 


MACRO OAI32xp5f_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI32xp5f_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.064 0.684 0.308 0.756 ; 
        RECT 0.064 0.108 0.252 0.18 ; 
        RECT 0.064 0.108 0.136 0.756 ; 
      LAYER M2 ; 
        RECT 0.152 0.684 0.672 0.756 ; 
      LAYER V1 ; 
        RECT 0.18 0.684 0.252 0.756 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.312 0.396 0.596 0.468 ; 
      LAYER M2 ; 
        RECT 0.244 0.396 0.652 0.468 ; 
      LAYER V1 ; 
        RECT 0.4 0.396 0.472 0.468 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.252 0.868 0.324 ; 
        RECT 0.532 0.54 0.792 0.612 ; 
        RECT 0.72 0.252 0.792 0.612 ; 
      LAYER M2 ; 
        RECT 0.588 0.252 0.996 0.324 ; 
      LAYER V1 ; 
        RECT 0.772 0.252 0.844 0.324 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.928 0.54 1.084 0.612 ; 
        RECT 0.928 0.392 1 0.612 ; 
      LAYER M2 ; 
        RECT 0.86 0.54 1.228 0.612 ; 
      LAYER V1 ; 
        RECT 0.996 0.54 1.068 0.612 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.236 0.396 1.308 0.584 ; 
        RECT 1.12 0.396 1.308 0.468 ; 
      LAYER M2 ; 
        RECT 0.972 0.396 1.38 0.468 ; 
      LAYER V1 ; 
        RECT 1.136 0.396 1.208 0.468 ; 
    END 
  END B2 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.684 1.452 0.756 ; 
        RECT 1.38 0.252 1.452 0.756 ; 
        RECT 1.044 0.252 1.452 0.324 ; 
        RECT 1.044 0.18 1.116 0.324 ; 
      LAYER M2 ; 
        RECT 0.836 0.684 1.352 0.756 ; 
      LAYER V1 ; 
        RECT 1.26 0.684 1.332 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.24 0.108 1.388 0.18 ; 
      RECT 0.376 0.108 0.92 0.18 ; 
    LAYER M2 ; 
      RECT 0.592 0.108 1.352 0.18 ; 
    LAYER V1 ; 
      RECT 1.26 0.108 1.332 0.18 ; 
      RECT 0.612 0.108 0.684 0.18 ; 
  END 
END OAI32xp5f_ASAP7_6t_SL 


MACRO OAI331xp33_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI331xp33_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.252 0.896 0.324 ; 
        RECT 0.72 0.252 0.792 0.584 ; 
      LAYER M2 ; 
        RECT 0.728 0.252 1.248 0.324 ; 
      LAYER V1 ; 
        RECT 0.8 0.252 0.872 0.324 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.62 0.756 ; 
        RECT 0.376 0.252 0.62 0.324 ; 
        RECT 0.504 0.252 0.576 0.756 ; 
      LAYER M2 ; 
        RECT 0.346 0.54 0.702 0.612 ; 
      LAYER V1 ; 
        RECT 0.504 0.54 0.576 0.612 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
      LAYER M2 ; 
        RECT 0.156 0.108 0.512 0.18 ; 
      LAYER V1 ; 
        RECT 0.18 0.108 0.252 0.18 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.396 1.084 0.468 ; 
        RECT 0.936 0.396 1.008 0.584 ; 
      LAYER M2 ; 
        RECT 0.612 0.396 1.244 0.468 ; 
      LAYER V1 ; 
        RECT 0.948 0.396 1.02 0.468 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.112 0.684 1.26 0.756 ; 
        RECT 1.152 0.512 1.224 0.756 ; 
      LAYER M2 ; 
        RECT 0.828 0.54 1.244 0.612 ; 
      LAYER V1 ; 
        RECT 1.152 0.54 1.224 0.612 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.684 1.516 0.756 ; 
        RECT 1.368 0.432 1.44 0.756 ; 
      LAYER M2 ; 
        RECT 1.368 0.54 1.68 0.612 ; 
      LAYER V1 ; 
        RECT 1.368 0.54 1.44 0.612 ; 
    END 
  END B3 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.648 0.304 1.72 0.584 ; 
      LAYER M2 ; 
        RECT 1.456 0.396 1.812 0.468 ; 
      LAYER V1 ; 
        RECT 1.648 0.396 1.72 0.468 ; 
    END 
  END C 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.64 0.684 1.872 0.756 ; 
        RECT 1.8 0.108 1.872 0.756 ; 
        RECT 1.672 0.108 1.872 0.18 ; 
        RECT 0.78 0.684 0.948 0.756 ; 
      LAYER M2 ; 
        RECT 0.804 0.684 1.788 0.756 ; 
      LAYER V1 ; 
        RECT 0.828 0.684 0.9 0.756 ; 
        RECT 1.692 0.684 1.764 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.044 0.252 1.548 0.324 ; 
      RECT 1.476 0.14 1.548 0.324 ; 
      RECT 0.396 0.108 1.332 0.18 ; 
  END 
END OAI331xp33_ASAP7_6t_SL 


MACRO OAI332xp33_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI332xp33_ASAP7_6t_SL 0 0 ; 
  SIZE 2.376 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.636 0.396 0.784 0.468 ; 
        RECT 0.376 0.684 0.708 0.756 ; 
        RECT 0.636 0.232 0.708 0.756 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.54 0.564 0.612 ; 
        RECT 0.492 0.252 0.564 0.612 ; 
        RECT 0.376 0.252 0.564 0.324 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.128 0.54 0.276 0.756 ; 
        RECT 0.204 0.108 0.276 0.756 ; 
        RECT 0.128 0.108 0.276 0.324 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.684 0.996 0.756 ; 
        RECT 0.924 0.252 0.996 0.756 ; 
        RECT 0.828 0.252 0.996 0.324 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.068 0.684 1.332 0.756 ; 
        RECT 1.068 0.396 1.288 0.468 ; 
        RECT 1.068 0.396 1.14 0.756 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.24 0.54 1.648 0.612 ; 
        RECT 1.428 0.396 1.648 0.468 ; 
        RECT 1.428 0.396 1.5 0.612 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.22 0.304 2.292 0.708 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.772 0.54 1.992 0.612 ; 
        RECT 1.92 0.396 1.992 0.612 ; 
        RECT 1.772 0.396 1.992 0.468 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.376 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.456 0.684 2.148 0.756 ; 
        RECT 2.076 0.252 2.148 0.756 ; 
        RECT 1.928 0.252 2.148 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.1 0.252 1.804 0.324 ; 
      RECT 1.732 0.108 1.804 0.324 ; 
      RECT 1.732 0.108 2.22 0.18 ; 
      RECT 0.804 0.108 1.568 0.18 ; 
      RECT 0.376 0.108 0.54 0.18 ; 
    LAYER M2 ; 
      RECT 0.376 0.108 0.936 0.18 ; 
    LAYER V1 ; 
      RECT 0.828 0.108 0.9 0.18 ; 
      RECT 0.396 0.108 0.468 0.18 ; 
  END 
END OAI332xp33_ASAP7_6t_SL 


MACRO OAI333xp33_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI333xp33_ASAP7_6t_SL 0 0 ; 
  SIZE 2.808 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.32 0.684 2.624 0.756 ; 
        RECT 2.552 0.348 2.624 0.756 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.236 0.54 2.468 0.612 ; 
        RECT 2.396 0.396 2.468 0.612 ; 
        RECT 2.236 0.396 2.468 0.468 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.792 0.396 2.088 0.468 ; 
        RECT 1.792 0.54 2.084 0.612 ; 
        RECT 1.792 0.396 1.864 0.612 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.684 1.02 0.756 ; 
        RECT 0.948 0.4 1.02 0.756 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.164 0.54 1.384 0.612 ; 
        RECT 1.312 0.396 1.384 0.612 ; 
        RECT 1.164 0.396 1.384 0.468 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.5 0.54 1.72 0.612 ; 
        RECT 1.648 0.396 1.72 0.612 ; 
        RECT 1.5 0.396 1.72 0.468 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.712 0.252 0.92 0.324 ; 
        RECT 0.636 0.512 0.784 0.596 ; 
        RECT 0.712 0.252 0.784 0.596 ; 
        RECT 0.376 0.684 0.708 0.756 ; 
        RECT 0.636 0.512 0.708 0.756 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.416 0.54 0.564 0.612 ; 
        RECT 0.492 0.252 0.564 0.612 ; 
        RECT 0.376 0.252 0.564 0.324 ; 
    END 
  END C2 
  PIN C3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.128 0.54 0.276 0.756 ; 
        RECT 0.204 0.108 0.276 0.756 ; 
        RECT 0.128 0.108 0.276 0.324 ; 
    END 
  END C3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.808 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.808 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 2.084 0.108 2.72 0.18 ; 
      LAYER M1 ; 
        RECT 2.696 0.108 2.768 0.652 ; 
        RECT 2.532 0.108 2.768 0.18 ; 
        RECT 2.02 0.108 2.216 0.18 ; 
      LAYER V1 ; 
        RECT 2.124 0.108 2.196 0.18 ; 
        RECT 2.556 0.108 2.628 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.06 0.252 2.412 0.324 ; 
      RECT 2.34 0.16 2.412 0.324 ; 
      RECT 1.06 0.16 1.132 0.324 ; 
      RECT 1.26 0.684 2.196 0.756 ; 
      RECT 1.26 0.108 1.572 0.18 ; 
      RECT 0.376 0.108 0.92 0.18 ; 
    LAYER M2 ; 
      RECT 0.808 0.108 1.572 0.18 ; 
    LAYER V1 ; 
      RECT 1.476 0.108 1.548 0.18 ; 
      RECT 0.828 0.108 0.9 0.18 ; 
  END 
END OAI333xp33_ASAP7_6t_SL 


MACRO OAI33xp5f_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI33xp5f_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.684 0.22 0.756 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.344 0.396 0.568 0.468 ; 
        RECT 0.344 0.684 0.492 0.756 ; 
        RECT 0.344 0.252 0.416 0.756 ; 
        RECT 0.26 0.252 0.416 0.324 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.536 0.54 0.792 0.612 ; 
        RECT 0.72 0.252 0.792 0.612 ; 
        RECT 0.644 0.252 0.792 0.324 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.008 0.684 1.248 0.756 ; 
        RECT 1.008 0.396 1.156 0.468 ; 
        RECT 1.008 0.396 1.08 0.756 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.376 0.684 1.524 0.756 ; 
        RECT 1.452 0.396 1.524 0.756 ; 
        RECT 1.284 0.396 1.524 0.468 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.76 0.684 1.908 0.756 ; 
        RECT 1.836 0.204 1.908 0.756 ; 
        RECT 1.648 0.396 1.908 0.468 ; 
    END 
  END B3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.864 0.252 1.764 0.324 ; 
        RECT 1.692 0.16 1.764 0.324 ; 
        RECT 0.704 0.684 0.936 0.756 ; 
        RECT 0.864 0.252 0.936 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.344 0.108 1.568 0.18 ; 
  END 
END OAI33xp5f_ASAP7_6t_SL 


MACRO OR2x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2x2_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.416 0.54 0.564 0.612 ; 
        RECT 0.492 0.252 0.564 0.612 ; 
        RECT 0.416 0.252 0.564 0.324 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.396 0.36 0.468 ; 
        RECT 0.072 0.684 0.272 0.756 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.684 1.224 0.756 ; 
        RECT 1.152 0.108 1.224 0.756 ; 
        RECT 0.808 0.108 1.224 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.396 0.684 0.708 0.756 ; 
      RECT 0.636 0.108 0.708 0.756 ; 
      RECT 0.636 0.396 0.904 0.468 ; 
      RECT 0.396 0.108 0.708 0.18 ; 
  END 
END OR2x2_ASAP7_6t_SL 


MACRO OR2x3R_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2x3R_ASAP7_6t_SL 0 0 ; 
  SIZE 2.592 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.612 0.252 0.684 0.44 ; 
        RECT 0.072 0.252 0.684 0.324 ; 
        RECT 0.072 0.684 0.276 0.756 ; 
        RECT 0.072 0.252 0.144 0.756 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.86 0.396 1.028 0.468 ; 
        RECT 0.376 0.54 0.936 0.612 ; 
        RECT 0.86 0.396 0.936 0.612 ; 
        RECT 0.376 0.54 0.524 0.756 ; 
        RECT 0.376 0.396 0.448 0.756 ; 
        RECT 0.288 0.396 0.448 0.468 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.592 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.26 0.684 2.52 0.756 ; 
        RECT 2.448 0.108 2.52 0.756 ; 
        RECT 1.148 0.108 2.52 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.808 0.684 1.136 0.756 ; 
      RECT 1.064 0.54 1.136 0.756 ; 
      RECT 1.064 0.54 1.224 0.612 ; 
      RECT 1.152 0.252 1.224 0.612 ; 
      RECT 0.936 0.252 1.224 0.324 ; 
      RECT 0.936 0.108 1.008 0.324 ; 
      RECT 0.376 0.108 1.008 0.18 ; 
  END 
END OR2x3R_ASAP7_6t_SL 


MACRO OR2x4_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2x4_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.464 0.576 0.612 ; 
        RECT 0.504 0.252 0.576 0.612 ; 
        RECT 0.376 0.252 0.576 0.324 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.464 0.304 0.612 ; 
        RECT 0.072 0.108 0.272 0.256 ; 
        RECT 0.072 0.108 0.144 0.612 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.828 0.684 1.656 0.756 ; 
        RECT 1.584 0.108 1.656 0.756 ; 
        RECT 0.828 0.108 1.656 0.18 ; 
        RECT 1.26 0.52 1.332 0.756 ; 
        RECT 1.26 0.108 1.332 0.344 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.684 0.72 0.756 ; 
      RECT 0.648 0.108 0.72 0.756 ; 
      RECT 0.648 0.396 0.792 0.468 ; 
      RECT 0.376 0.108 0.72 0.18 ; 
  END 
END OR2x4_ASAP7_6t_SL 


MACRO OR3x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR3x1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.296 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.252 0.22 0.324 ; 
        RECT 0.072 0.252 0.144 0.756 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.396 0.576 0.468 ; 
        RECT 0.352 0.608 0.5 0.756 ; 
        RECT 0.428 0.252 0.5 0.756 ; 
        RECT 0.352 0.252 0.5 0.324 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.644 0.54 0.792 0.612 ; 
        RECT 0.72 0.252 0.792 0.612 ; 
        RECT 0.644 0.252 0.792 0.324 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.296 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.044 0.684 1.224 0.756 ; 
        RECT 1.152 0.108 1.224 0.756 ; 
        RECT 1.044 0.108 1.224 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.612 0.684 0.936 0.756 ; 
      RECT 0.864 0.108 0.936 0.756 ; 
      RECT 0.864 0.396 1.048 0.468 ; 
      RECT 0.16 0.108 0.936 0.18 ; 
  END 
END OR3x1_ASAP7_6t_SL 


MACRO OR3x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR3x2_ASAP7_6t_SL 0 0 ; 
  SIZE 1.512 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.252 0.22 0.324 ; 
        RECT 0.072 0.252 0.144 0.756 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.42 0.396 0.572 0.468 ; 
        RECT 0.344 0.608 0.492 0.756 ; 
        RECT 0.42 0.252 0.492 0.756 ; 
        RECT 0.344 0.252 0.492 0.324 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.632 0.54 0.78 0.612 ; 
        RECT 0.708 0.252 0.78 0.612 ; 
        RECT 0.632 0.252 0.78 0.324 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.512 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.684 1.44 0.756 ; 
        RECT 1.368 0.108 1.44 0.756 ; 
        RECT 1.024 0.108 1.44 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.592 0.684 0.924 0.756 ; 
      RECT 0.852 0.108 0.924 0.756 ; 
      RECT 0.852 0.396 1.136 0.468 ; 
      RECT 0.16 0.108 0.924 0.18 ; 
  END 
END OR3x2_ASAP7_6t_SL 


MACRO OR3x4_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR3x4_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.608 0.272 0.756 ; 
        RECT 0.072 0.252 0.272 0.4 ; 
        RECT 0.072 0.252 0.144 0.756 ; 
      LAYER M2 ; 
        RECT 0.072 0.252 0.356 0.324 ; 
      LAYER V1 ; 
        RECT 0.156 0.252 0.228 0.324 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.356 0.412 0.584 0.484 ; 
        RECT 0.356 0.412 0.504 0.756 ; 
      LAYER M2 ; 
        RECT 0.268 0.54 0.688 0.612 ; 
      LAYER V1 ; 
        RECT 0.384 0.54 0.456 0.612 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.252 0.792 0.488 ; 
        RECT 0.376 0.252 0.792 0.324 ; 
      LAYER M2 ; 
        RECT 0.6 0.396 0.896 0.468 ; 
      LAYER V1 ; 
        RECT 0.72 0.396 0.792 0.468 ; 
    END 
  END C 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.044 0.684 1.872 0.756 ; 
        RECT 1.8 0.108 1.872 0.756 ; 
        RECT 1.044 0.108 1.872 0.18 ; 
        RECT 1.476 0.52 1.548 0.756 ; 
        RECT 1.476 0.108 1.548 0.344 ; 
      LAYER M2 ; 
        RECT 1.392 0.396 1.872 0.468 ; 
      LAYER V1 ; 
        RECT 1.8 0.396 1.872 0.468 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.612 0.684 0.936 0.756 ; 
      RECT 0.864 0.108 0.936 0.756 ; 
      RECT 0.864 0.396 1.012 0.468 ; 
      RECT 0.16 0.108 0.936 0.18 ; 
  END 
END OR3x4_ASAP7_6t_SL 


MACRO OR4x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR4x1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.036 0.604 0.252 0.752 ; 
        RECT 0.036 0.108 0.252 0.256 ; 
        RECT 0.036 0.396 0.188 0.468 ; 
        RECT 0.036 0.108 0.108 0.752 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.324 0.396 0.576 0.468 ; 
        RECT 0.324 0.608 0.472 0.756 ; 
        RECT 0.324 0.252 0.472 0.468 ; 
        RECT 0.324 0.252 0.396 0.756 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.544 0.54 0.792 0.612 ; 
        RECT 0.72 0.252 0.792 0.612 ; 
        RECT 0.64 0.252 0.792 0.324 ; 
        RECT 0.544 0.54 0.692 0.756 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.908 0.54 1.056 0.612 ; 
        RECT 0.908 0.252 1.056 0.324 ; 
        RECT 0.94 0.252 1.012 0.612 ; 
    END 
  END D 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.3 0.684 1.568 0.756 ; 
        RECT 1.3 0.108 1.568 0.18 ; 
        RECT 1.3 0.108 1.372 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.828 0.684 1.228 0.756 ; 
      RECT 1.156 0.108 1.228 0.756 ; 
      RECT 0.376 0.108 1.228 0.18 ; 
  END 
END OR4x1_ASAP7_6t_SL 


MACRO OR4x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR4x2_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.544 0.68 1.692 0.752 ; 
        RECT 1.62 0.108 1.692 0.752 ; 
        RECT 1.54 0.396 1.692 0.468 ; 
        RECT 1.456 0.108 1.692 0.18 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.244 0.608 1.44 0.756 ; 
        RECT 1.368 0.324 1.44 0.756 ; 
        RECT 1.272 0.252 1.42 0.468 ; 
        RECT 1.152 0.396 1.44 0.468 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.54 1.172 0.756 ; 
        RECT 0.936 0.252 1.088 0.324 ; 
        RECT 0.936 0.54 1.172 0.612 ; 
        RECT 0.936 0.252 1.008 0.612 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.664 0.54 0.812 0.612 ; 
        RECT 0.664 0.252 0.812 0.324 ; 
        RECT 0.716 0.252 0.788 0.612 ; 
    END 
  END D 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.16 0.684 0.42 0.756 ; 
        RECT 0.348 0.108 0.42 0.756 ; 
        RECT 0.16 0.108 0.42 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.492 0.684 0.9 0.756 ; 
      RECT 0.492 0.108 0.564 0.756 ; 
      RECT 0.492 0.108 1.332 0.18 ; 
  END 
END OR4x2_ASAP7_6t_SL 


MACRO OR5x1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR5x1_ASAP7_6t_SL 0 0 ; 
  SIZE 1.728 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.064 0.684 0.26 0.756 ; 
        RECT 0.064 0.172 0.136 0.756 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.388 0.684 0.564 0.756 ; 
        RECT 0.492 0.252 0.564 0.756 ; 
        RECT 0.412 0.252 0.564 0.324 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.712 0.684 0.908 0.756 ; 
        RECT 0.712 0.252 0.784 0.756 ; 
        RECT 0.636 0.252 0.784 0.4 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.008 0.656 1.156 0.756 ; 
        RECT 1.008 0.528 1.08 0.756 ; 
        RECT 0.924 0.528 1.08 0.6 ; 
        RECT 0.856 0.252 1.004 0.4 ; 
        RECT 0.924 0.252 0.996 0.6 ; 
    END 
  END D 
  PIN E 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.284 0.504 1.356 0.728 ; 
        RECT 1.18 0.252 1.336 0.324 ; 
        RECT 1.18 0.504 1.356 0.576 ; 
        RECT 1.18 0.252 1.252 0.576 ; 
    END 
  END E 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.728 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.468 0.684 1.664 0.756 ; 
        RECT 1.592 0.208 1.664 0.756 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.284 0.428 0.356 0.6 ; 
      RECT 0.208 0.428 0.356 0.5 ; 
      RECT 1.436 0.108 1.508 0.456 ; 
      RECT 0.208 0.108 0.28 0.5 ; 
      RECT 0.208 0.108 1.508 0.18 ; 
  END 
END OR5x1_ASAP7_6t_SL 


MACRO OR5x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR5x2_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.144 0.604 0.292 0.752 ; 
        RECT 0.144 0.252 0.292 0.4 ; 
        RECT 0.144 0.252 0.216 0.752 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.604 0.572 0.752 ; 
        RECT 0.5 0.252 0.572 0.752 ; 
        RECT 0.376 0.252 0.572 0.4 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.604 0.92 0.752 ; 
        RECT 0.72 0.448 0.792 0.752 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.928 0.252 1 0.464 ; 
        RECT 0.808 0.252 1 0.324 ; 
    END 
  END D 
  PIN E 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.032 0.54 1.276 0.612 ; 
        RECT 1.152 0.396 1.224 0.612 ; 
    END 
  END E 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.524 0.684 1.872 0.756 ; 
        RECT 1.8 0.108 1.872 0.756 ; 
        RECT 1.524 0.108 1.872 0.18 ; 
        RECT 1.524 0.536 1.596 0.756 ; 
        RECT 1.524 0.108 1.596 0.328 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.024 0.684 1.448 0.756 ; 
      RECT 1.376 0.108 1.448 0.756 ; 
      RECT 0.132 0.108 1.448 0.18 ; 
  END 
END OR5x2_ASAP7_6t_SL 


MACRO SDFHx1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN SDFHx1_ASAP7_6t_SL 0 0 ; 
  SIZE 5.832 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 1.044 0.684 1.2 0.756 ; 
        RECT 1.044 0.54 1.116 0.756 ; 
        RECT 0.936 0.108 1.084 0.184 ; 
        RECT 0.936 0.54 1.116 0.612 ; 
        RECT 0.936 0.108 1.008 0.612 ; 
      LAYER M2 ; 
        RECT 0.54 0.54 1.432 0.612 ; 
      LAYER V1 ; 
        RECT 0.988 0.54 1.06 0.612 ; 
    END 
  END CLK 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.56 0.684 5.76 0.756 ; 
        RECT 5.688 0.108 5.76 0.756 ; 
        RECT 5.5 0.108 5.76 0.18 ; 
    END 
  END QN 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.48 0.396 1.656 0.468 ; 
        RECT 1.48 0.108 1.564 0.468 ; 
        RECT 1.308 0.108 1.564 0.18 ; 
        RECT 0.072 0.108 0.276 0.18 ; 
        RECT 0.072 0.684 0.22 0.756 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
      LAYER M2 ; 
        RECT 0.08 0.108 1.592 0.18 ; 
      LAYER V1 ; 
        RECT 0.18 0.108 0.252 0.18 ; 
        RECT 1.476 0.108 1.548 0.18 ; 
    END 
  END SE 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 5.832 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.832 0.036 ; 
    END 
  END VSS 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.212 0.396 2.416 0.468 ; 
      LAYER M2 ; 
        RECT 2.008 0.396 2.528 0.468 ; 
      LAYER V1 ; 
        RECT 2.268 0.396 2.34 0.468 ; 
    END 
  END D 
  PIN SI 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.716 0.396 2.788 0.66 ; 
        RECT 2.548 0.396 2.788 0.468 ; 
      LAYER M2 ; 
        RECT 2.652 0.396 3.172 0.468 ; 
      LAYER V1 ; 
        RECT 2.692 0.396 2.764 0.468 ; 
    END 
  END SI 
  OBS 
    LAYER M1 ; 
      RECT 5.472 0.252 5.544 0.5 ; 
      RECT 5.416 0.252 5.564 0.324 ; 
      RECT 4.912 0.684 5.272 0.756 ; 
      RECT 5.2 0.108 5.272 0.756 ; 
      RECT 4.608 0.28 4.8 0.352 ; 
      RECT 4.728 0.108 4.8 0.352 ; 
      RECT 4.728 0.108 5.272 0.18 ; 
      RECT 5.036 0.252 5.108 0.504 ; 
      RECT 4.932 0.252 5.108 0.324 ; 
      RECT 4.264 0.68 4.464 0.752 ; 
      RECT 4.392 0.108 4.464 0.752 ; 
      RECT 4.048 0.108 4.464 0.18 ; 
      RECT 4.176 0.252 4.248 0.492 ; 
      RECT 4.128 0.252 4.288 0.324 ; 
      RECT 3.916 0.54 4.072 0.612 ; 
      RECT 3.96 0.376 4.032 0.612 ; 
      RECT 3.6 0.684 4.024 0.756 ; 
      RECT 3.6 0.188 3.672 0.756 ; 
      RECT 3.488 0.308 3.672 0.38 ; 
      RECT 3.6 0.188 3.924 0.26 ; 
      RECT 2.94 0.684 3.368 0.756 ; 
      RECT 3.296 0.108 3.368 0.756 ; 
      RECT 3.204 0.108 3.368 0.18 ; 
      RECT 3.096 0.252 3.168 0.464 ; 
      RECT 3.048 0.252 3.168 0.324 ; 
      RECT 2.888 0.54 3.036 0.612 ; 
      RECT 2.888 0.392 2.96 0.612 ; 
      RECT 2.264 0.252 2.832 0.324 ; 
      RECT 2.76 0.16 2.832 0.324 ; 
      RECT 2.76 0.16 2.948 0.232 ; 
      RECT 1.692 0.684 2.644 0.756 ; 
      RECT 2.572 0.592 2.644 0.756 ; 
      RECT 1.328 0.684 1.548 0.756 ; 
      RECT 1.328 0.54 1.4 0.756 ; 
      RECT 1.328 0.54 1.736 0.612 ; 
      RECT 1.156 0.396 1.38 0.468 ; 
      RECT 1.308 0.252 1.38 0.468 ; 
      RECT 1.156 0.252 1.38 0.324 ; 
      RECT 0.612 0.684 0.776 0.756 ; 
      RECT 0.704 0.108 0.776 0.756 ; 
      RECT 0.612 0.108 0.776 0.18 ; 
      RECT 0.324 0.684 0.488 0.756 ; 
      RECT 0.324 0.252 0.396 0.756 ; 
      RECT 0.324 0.252 0.488 0.324 ; 
      RECT 4.608 0.452 4.68 0.688 ; 
      RECT 3.744 0.38 3.816 0.576 ; 
      RECT 3.456 0.504 3.528 0.688 ; 
      RECT 1.692 0.108 2.628 0.18 ; 
      RECT 1.86 0.54 2.448 0.612 ; 
      RECT 1.78 0.396 2.088 0.468 ; 
    LAYER M2 ; 
      RECT 4.392 0.252 5.564 0.324 ; 
      RECT 1.584 0.54 4.68 0.612 ; 
      RECT 0.612 0.252 4.248 0.324 ; 
      RECT 3.296 0.396 3.816 0.468 ; 
      RECT 0.292 0.396 1.88 0.468 ; 
    LAYER V1 ; 
      RECT 5.472 0.252 5.544 0.324 ; 
      RECT 5.016 0.252 5.088 0.324 ; 
      RECT 4.608 0.54 4.68 0.612 ; 
      RECT 4.392 0.252 4.464 0.324 ; 
      RECT 4.176 0.252 4.248 0.324 ; 
      RECT 3.96 0.54 4.032 0.612 ; 
      RECT 3.744 0.396 3.816 0.468 ; 
      RECT 3.456 0.54 3.528 0.612 ; 
      RECT 3.296 0.396 3.368 0.468 ; 
      RECT 3.076 0.252 3.148 0.324 ; 
      RECT 2.912 0.54 2.984 0.612 ; 
      RECT 1.808 0.396 1.88 0.468 ; 
      RECT 1.584 0.54 1.656 0.612 ; 
      RECT 1.264 0.252 1.336 0.324 ; 
      RECT 0.704 0.252 0.776 0.324 ; 
      RECT 0.324 0.396 0.396 0.468 ; 
  END 
END SDFHx1_ASAP7_6t_SL 


MACRO SDFHx2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN SDFHx2_ASAP7_6t_SL 0 0 ; 
  SIZE 6.048 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 4.824 0.684 5.304 0.756 ; 
        RECT 5.232 0.108 5.304 0.756 ; 
        RECT 5.128 0.108 5.304 0.184 ; 
        RECT 4.824 0.376 4.896 0.756 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.32 0.396 1.54 0.468 ; 
        RECT 1.32 0.248 1.392 0.468 ; 
        RECT 1.148 0.248 1.392 0.324 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.56 0.684 5.76 0.756 ; 
        RECT 5.688 0.108 5.76 0.756 ; 
        RECT 5.5 0.108 5.76 0.18 ; 
    END 
  END QN 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.396 0.74 0.468 ; 
        RECT 0.128 0.684 0.664 0.756 ; 
        RECT 0.592 0.396 0.664 0.756 ; 
        RECT 0.128 0.108 0.276 0.18 ; 
        RECT 0.128 0.108 0.2 0.756 ; 
    END 
  END SE 
  PIN SI 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.672 0.684 1.936 0.756 ; 
        RECT 1.864 0.396 1.936 0.756 ; 
        RECT 1.672 0.396 1.936 0.468 ; 
    END 
  END SI 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 6.048 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 6.048 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 4.968 0.54 5.132 0.612 ; 
      RECT 4.968 0.204 5.04 0.612 ; 
      RECT 4.608 0.204 4.68 0.488 ; 
      RECT 4.608 0.204 5.04 0.276 ; 
      RECT 3.888 0.684 4.16 0.756 ; 
      RECT 3.888 0.108 3.96 0.756 ; 
      RECT 3.74 0.28 3.96 0.352 ; 
      RECT 3.888 0.108 4.16 0.18 ; 
      RECT 3.4 0.68 3.64 0.752 ; 
      RECT 3.568 0.108 3.64 0.752 ; 
      RECT 3.184 0.108 3.64 0.18 ; 
      RECT 3.312 0.252 3.384 0.492 ; 
      RECT 3.264 0.252 3.424 0.324 ; 
      RECT 3.052 0.54 3.208 0.612 ; 
      RECT 3.096 0.376 3.168 0.612 ; 
      RECT 2.736 0.684 3.16 0.756 ; 
      RECT 2.736 0.188 2.808 0.756 ; 
      RECT 2.664 0.308 2.808 0.38 ; 
      RECT 2.736 0.188 3.06 0.26 ; 
      RECT 2.124 0.684 2.504 0.756 ; 
      RECT 2.432 0.108 2.504 0.756 ; 
      RECT 2.34 0.108 2.504 0.18 ; 
      RECT 2.224 0.252 2.296 0.464 ; 
      RECT 2.148 0.252 2.296 0.324 ; 
      RECT 1.464 0.252 2.004 0.324 ; 
      RECT 1.932 0.108 2.004 0.324 ; 
      RECT 1.464 0.16 1.536 0.324 ; 
      RECT 1.932 0.108 2.196 0.18 ; 
      RECT 2.028 0.54 2.176 0.612 ; 
      RECT 2.028 0.408 2.1 0.612 ; 
      RECT 0.828 0.54 0.9 0.712 ; 
      RECT 0.828 0.54 1.764 0.612 ; 
      RECT 0.344 0.54 0.492 0.612 ; 
      RECT 0.344 0.252 0.42 0.612 ; 
      RECT 0.912 0.396 1.196 0.468 ; 
      RECT 0.912 0.252 0.984 0.468 ; 
      RECT 0.344 0.252 0.984 0.324 ; 
      RECT 5.472 0.352 5.544 0.5 ; 
      RECT 4.464 0.232 4.536 0.632 ; 
      RECT 4.032 0.356 4.104 0.504 ; 
      RECT 3.74 0.452 3.812 0.688 ; 
      RECT 2.88 0.38 2.952 0.576 ; 
      RECT 2.592 0.504 2.664 0.688 ; 
      RECT 1.66 0.108 1.808 0.18 ; 
      RECT 1.044 0.684 1.548 0.756 ; 
      RECT 0.792 0.108 0.94 0.18 ; 
    LAYER M2 ; 
      RECT 3.548 0.396 5.564 0.468 ; 
      RECT 2.18 0.252 4.7 0.324 ; 
      RECT 2.048 0.54 4.556 0.612 ; 
      RECT 2.432 0.396 2.952 0.468 ; 
      RECT 0.768 0.108 1.86 0.18 ; 
    LAYER V1 ; 
      RECT 5.472 0.396 5.544 0.468 ; 
      RECT 4.608 0.252 4.68 0.324 ; 
      RECT 4.464 0.54 4.536 0.612 ; 
      RECT 4.032 0.396 4.104 0.468 ; 
      RECT 3.74 0.54 3.812 0.612 ; 
      RECT 3.568 0.396 3.64 0.468 ; 
      RECT 3.312 0.252 3.384 0.324 ; 
      RECT 3.096 0.54 3.168 0.612 ; 
      RECT 2.88 0.396 2.952 0.468 ; 
      RECT 2.592 0.54 2.664 0.612 ; 
      RECT 2.432 0.396 2.504 0.468 ; 
      RECT 2.2 0.252 2.272 0.324 ; 
      RECT 2.068 0.54 2.14 0.612 ; 
      RECT 1.692 0.108 1.764 0.18 ; 
      RECT 0.828 0.108 0.9 0.18 ; 
  END 
END SDFHx2_ASAP7_6t_SL 


MACRO SDFHx3_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN SDFHx3_ASAP7_6t_SL 0 0 ; 
  SIZE 6.264 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 4.824 0.684 5.304 0.756 ; 
        RECT 5.232 0.108 5.304 0.756 ; 
        RECT 5.128 0.108 5.304 0.184 ; 
        RECT 4.824 0.376 4.896 0.756 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.32 0.396 1.54 0.468 ; 
        RECT 1.32 0.248 1.392 0.468 ; 
        RECT 1.148 0.248 1.392 0.324 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.56 0.684 6.192 0.756 ; 
        RECT 6.12 0.108 6.192 0.756 ; 
        RECT 5.5 0.108 6.192 0.18 ; 
    END 
  END QN 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.396 0.74 0.468 ; 
        RECT 0.128 0.684 0.664 0.756 ; 
        RECT 0.592 0.396 0.664 0.756 ; 
        RECT 0.128 0.108 0.276 0.18 ; 
        RECT 0.128 0.108 0.2 0.756 ; 
    END 
  END SE 
  PIN SI 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.672 0.684 1.936 0.756 ; 
        RECT 1.864 0.396 1.936 0.756 ; 
        RECT 1.672 0.396 1.936 0.468 ; 
    END 
  END SI 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 6.264 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 6.264 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 4.968 0.54 5.132 0.612 ; 
      RECT 4.968 0.204 5.04 0.612 ; 
      RECT 4.608 0.204 4.68 0.488 ; 
      RECT 4.608 0.204 5.04 0.276 ; 
      RECT 3.888 0.684 4.16 0.756 ; 
      RECT 3.888 0.108 3.96 0.756 ; 
      RECT 3.74 0.28 3.96 0.352 ; 
      RECT 3.888 0.108 4.16 0.18 ; 
      RECT 3.4 0.68 3.64 0.752 ; 
      RECT 3.568 0.108 3.64 0.752 ; 
      RECT 3.184 0.108 3.64 0.18 ; 
      RECT 3.312 0.252 3.384 0.492 ; 
      RECT 3.264 0.252 3.424 0.324 ; 
      RECT 3.052 0.54 3.208 0.612 ; 
      RECT 3.096 0.376 3.168 0.612 ; 
      RECT 2.736 0.684 3.16 0.756 ; 
      RECT 2.736 0.188 2.808 0.756 ; 
      RECT 2.664 0.308 2.808 0.38 ; 
      RECT 2.736 0.188 3.06 0.26 ; 
      RECT 2.124 0.684 2.504 0.756 ; 
      RECT 2.432 0.108 2.504 0.756 ; 
      RECT 2.34 0.108 2.504 0.18 ; 
      RECT 2.224 0.252 2.296 0.464 ; 
      RECT 2.148 0.252 2.296 0.324 ; 
      RECT 1.464 0.252 2.004 0.324 ; 
      RECT 1.932 0.108 2.004 0.324 ; 
      RECT 1.464 0.16 1.536 0.324 ; 
      RECT 1.932 0.108 2.196 0.18 ; 
      RECT 2.028 0.54 2.176 0.612 ; 
      RECT 2.028 0.408 2.1 0.612 ; 
      RECT 0.828 0.54 0.9 0.712 ; 
      RECT 0.828 0.54 1.764 0.612 ; 
      RECT 0.344 0.54 0.492 0.612 ; 
      RECT 0.344 0.252 0.42 0.612 ; 
      RECT 0.912 0.396 1.196 0.468 ; 
      RECT 0.912 0.252 0.984 0.468 ; 
      RECT 0.344 0.252 0.984 0.324 ; 
      RECT 5.432 0.396 6.008 0.468 ; 
      RECT 4.464 0.232 4.536 0.632 ; 
      RECT 4.032 0.356 4.104 0.504 ; 
      RECT 3.74 0.452 3.812 0.688 ; 
      RECT 2.88 0.38 2.952 0.576 ; 
      RECT 2.592 0.504 2.664 0.688 ; 
      RECT 1.66 0.108 1.808 0.18 ; 
      RECT 1.044 0.684 1.548 0.756 ; 
      RECT 0.792 0.108 0.94 0.18 ; 
    LAYER M2 ; 
      RECT 3.548 0.396 5.564 0.468 ; 
      RECT 2.18 0.252 4.7 0.324 ; 
      RECT 2.048 0.54 4.556 0.612 ; 
      RECT 2.432 0.396 2.952 0.468 ; 
      RECT 0.768 0.108 1.86 0.18 ; 
    LAYER V1 ; 
      RECT 5.472 0.396 5.544 0.468 ; 
      RECT 4.608 0.252 4.68 0.324 ; 
      RECT 4.464 0.54 4.536 0.612 ; 
      RECT 4.032 0.396 4.104 0.468 ; 
      RECT 3.74 0.54 3.812 0.612 ; 
      RECT 3.568 0.396 3.64 0.468 ; 
      RECT 3.312 0.252 3.384 0.324 ; 
      RECT 3.096 0.54 3.168 0.612 ; 
      RECT 2.88 0.396 2.952 0.468 ; 
      RECT 2.592 0.54 2.664 0.612 ; 
      RECT 2.432 0.396 2.504 0.468 ; 
      RECT 2.2 0.252 2.272 0.324 ; 
      RECT 2.068 0.54 2.14 0.612 ; 
      RECT 1.692 0.108 1.764 0.18 ; 
      RECT 0.828 0.108 0.9 0.18 ; 
  END 
END SDFHx3_ASAP7_6t_SL 


MACRO SDFHx4_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN SDFHx4_ASAP7_6t_SL 0 0 ; 
  SIZE 6.48 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 4.824 0.684 5.304 0.756 ; 
        RECT 5.232 0.108 5.304 0.756 ; 
        RECT 5.128 0.108 5.304 0.184 ; 
        RECT 4.824 0.376 4.896 0.756 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.32 0.396 1.54 0.468 ; 
        RECT 1.32 0.248 1.392 0.468 ; 
        RECT 1.148 0.248 1.392 0.324 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.56 0.684 6.304 0.756 ; 
        RECT 6.232 0.108 6.304 0.756 ; 
        RECT 5.56 0.108 6.304 0.18 ; 
    END 
  END QN 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.396 0.74 0.468 ; 
        RECT 0.128 0.684 0.664 0.756 ; 
        RECT 0.592 0.396 0.664 0.756 ; 
        RECT 0.128 0.108 0.276 0.18 ; 
        RECT 0.128 0.108 0.2 0.756 ; 
    END 
  END SE 
  PIN SI 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.672 0.684 1.936 0.756 ; 
        RECT 1.864 0.396 1.936 0.756 ; 
        RECT 1.672 0.396 1.936 0.468 ; 
    END 
  END SI 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 6.48 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 6.48 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 4.968 0.54 5.132 0.612 ; 
      RECT 4.968 0.204 5.04 0.612 ; 
      RECT 4.608 0.204 4.68 0.488 ; 
      RECT 4.608 0.204 5.04 0.276 ; 
      RECT 3.888 0.684 4.16 0.756 ; 
      RECT 3.888 0.108 3.96 0.756 ; 
      RECT 3.74 0.28 3.96 0.352 ; 
      RECT 3.888 0.108 4.16 0.18 ; 
      RECT 3.4 0.68 3.64 0.752 ; 
      RECT 3.568 0.108 3.64 0.752 ; 
      RECT 3.184 0.108 3.64 0.18 ; 
      RECT 3.312 0.252 3.384 0.492 ; 
      RECT 3.264 0.252 3.424 0.324 ; 
      RECT 3.052 0.54 3.208 0.612 ; 
      RECT 3.096 0.376 3.168 0.612 ; 
      RECT 2.736 0.684 3.16 0.756 ; 
      RECT 2.736 0.188 2.808 0.756 ; 
      RECT 2.664 0.308 2.808 0.38 ; 
      RECT 2.736 0.188 3.06 0.26 ; 
      RECT 2.124 0.684 2.504 0.756 ; 
      RECT 2.432 0.108 2.504 0.756 ; 
      RECT 2.34 0.108 2.504 0.18 ; 
      RECT 2.224 0.252 2.296 0.464 ; 
      RECT 2.148 0.252 2.296 0.324 ; 
      RECT 1.464 0.252 2.004 0.324 ; 
      RECT 1.932 0.108 2.004 0.324 ; 
      RECT 1.464 0.16 1.536 0.324 ; 
      RECT 1.932 0.108 2.196 0.18 ; 
      RECT 2.028 0.54 2.176 0.612 ; 
      RECT 2.028 0.408 2.1 0.612 ; 
      RECT 0.828 0.54 0.9 0.712 ; 
      RECT 0.828 0.54 1.764 0.612 ; 
      RECT 0.344 0.54 0.492 0.612 ; 
      RECT 0.344 0.252 0.42 0.612 ; 
      RECT 0.912 0.396 1.196 0.468 ; 
      RECT 0.912 0.252 0.984 0.468 ; 
      RECT 0.344 0.252 0.984 0.324 ; 
      RECT 5.452 0.396 6.104 0.468 ; 
      RECT 4.464 0.232 4.536 0.632 ; 
      RECT 4.032 0.356 4.104 0.504 ; 
      RECT 3.74 0.452 3.812 0.688 ; 
      RECT 2.88 0.38 2.952 0.576 ; 
      RECT 2.592 0.504 2.664 0.688 ; 
      RECT 1.66 0.108 1.808 0.18 ; 
      RECT 1.044 0.684 1.548 0.756 ; 
      RECT 0.792 0.108 0.94 0.18 ; 
    LAYER M2 ; 
      RECT 3.548 0.396 5.564 0.468 ; 
      RECT 2.18 0.252 4.7 0.324 ; 
      RECT 2.048 0.54 4.556 0.612 ; 
      RECT 2.432 0.396 2.952 0.468 ; 
      RECT 0.768 0.108 1.86 0.18 ; 
    LAYER V1 ; 
      RECT 5.472 0.396 5.544 0.468 ; 
      RECT 4.608 0.252 4.68 0.324 ; 
      RECT 4.464 0.54 4.536 0.612 ; 
      RECT 4.032 0.396 4.104 0.468 ; 
      RECT 3.74 0.54 3.812 0.612 ; 
      RECT 3.568 0.396 3.64 0.468 ; 
      RECT 3.312 0.252 3.384 0.324 ; 
      RECT 3.096 0.54 3.168 0.612 ; 
      RECT 2.88 0.396 2.952 0.468 ; 
      RECT 2.592 0.54 2.664 0.612 ; 
      RECT 2.432 0.396 2.504 0.468 ; 
      RECT 2.2 0.252 2.272 0.324 ; 
      RECT 2.068 0.54 2.14 0.612 ; 
      RECT 1.692 0.108 1.764 0.18 ; 
      RECT 0.828 0.108 0.9 0.18 ; 
  END 
END SDFHx4_ASAP7_6t_SL 


MACRO SDFLx1_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN SDFLx1_ASAP7_6t_SL 0 0 ; 
  SIZE 5.832 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 4.824 0.684 5.304 0.756 ; 
        RECT 5.232 0.108 5.304 0.756 ; 
        RECT 5.128 0.108 5.304 0.184 ; 
        RECT 4.824 0.376 4.896 0.756 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.32 0.396 1.54 0.468 ; 
        RECT 1.32 0.248 1.392 0.468 ; 
        RECT 1.148 0.248 1.392 0.324 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.56 0.684 5.76 0.756 ; 
        RECT 5.688 0.108 5.76 0.756 ; 
        RECT 5.54 0.108 5.76 0.18 ; 
    END 
  END QN 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.396 0.74 0.468 ; 
        RECT 0.128 0.684 0.664 0.756 ; 
        RECT 0.592 0.396 0.664 0.756 ; 
        RECT 0.128 0.108 0.276 0.18 ; 
        RECT 0.128 0.108 0.2 0.756 ; 
    END 
  END SE 
  PIN SI 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.672 0.684 1.936 0.756 ; 
        RECT 1.864 0.396 1.936 0.756 ; 
        RECT 1.672 0.396 1.936 0.468 ; 
    END 
  END SI 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 5.832 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.832 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 4.608 0.204 4.68 0.632 ; 
      RECT 4.968 0.54 5.132 0.612 ; 
      RECT 4.968 0.204 5.04 0.612 ; 
      RECT 4.608 0.204 5.04 0.276 ; 
      RECT 3.888 0.684 4.16 0.756 ; 
      RECT 3.888 0.108 3.96 0.756 ; 
      RECT 3.74 0.28 3.96 0.352 ; 
      RECT 3.888 0.108 4.16 0.18 ; 
      RECT 3.4 0.68 3.64 0.752 ; 
      RECT 3.568 0.108 3.64 0.752 ; 
      RECT 3.184 0.108 3.64 0.18 ; 
      RECT 3.312 0.252 3.384 0.492 ; 
      RECT 3.264 0.252 3.424 0.324 ; 
      RECT 3.052 0.54 3.208 0.612 ; 
      RECT 3.096 0.376 3.168 0.612 ; 
      RECT 2.736 0.684 3.16 0.756 ; 
      RECT 2.736 0.188 2.808 0.756 ; 
      RECT 2.664 0.308 2.808 0.38 ; 
      RECT 2.736 0.188 3.06 0.26 ; 
      RECT 2.124 0.684 2.504 0.756 ; 
      RECT 2.432 0.108 2.504 0.756 ; 
      RECT 2.34 0.108 2.504 0.18 ; 
      RECT 2.224 0.252 2.296 0.464 ; 
      RECT 2.148 0.252 2.296 0.324 ; 
      RECT 1.464 0.252 2.004 0.324 ; 
      RECT 1.932 0.108 2.004 0.324 ; 
      RECT 1.464 0.16 1.536 0.324 ; 
      RECT 1.932 0.108 2.196 0.18 ; 
      RECT 2.028 0.54 2.176 0.612 ; 
      RECT 2.028 0.408 2.1 0.612 ; 
      RECT 0.828 0.54 0.9 0.712 ; 
      RECT 0.828 0.54 1.764 0.612 ; 
      RECT 0.344 0.54 0.492 0.612 ; 
      RECT 0.344 0.252 0.42 0.612 ; 
      RECT 0.912 0.396 1.196 0.468 ; 
      RECT 0.912 0.252 0.984 0.468 ; 
      RECT 0.344 0.252 0.984 0.324 ; 
      RECT 5.472 0.352 5.544 0.5 ; 
      RECT 4.464 0.232 4.536 0.632 ; 
      RECT 4.032 0.356 4.104 0.504 ; 
      RECT 3.74 0.452 3.812 0.688 ; 
      RECT 2.88 0.38 2.952 0.576 ; 
      RECT 2.592 0.504 2.664 0.688 ; 
      RECT 1.66 0.108 1.808 0.18 ; 
      RECT 1.044 0.684 1.548 0.756 ; 
      RECT 0.792 0.108 0.94 0.18 ; 
    LAYER M2 ; 
      RECT 3.548 0.396 5.564 0.468 ; 
      RECT 2.048 0.54 4.7 0.612 ; 
      RECT 2.18 0.252 4.556 0.324 ; 
      RECT 2.432 0.396 2.952 0.468 ; 
      RECT 0.768 0.108 1.86 0.18 ; 
    LAYER V1 ; 
      RECT 5.472 0.396 5.544 0.468 ; 
      RECT 4.608 0.54 4.68 0.612 ; 
      RECT 4.464 0.252 4.536 0.324 ; 
      RECT 4.032 0.396 4.104 0.468 ; 
      RECT 3.74 0.54 3.812 0.612 ; 
      RECT 3.568 0.396 3.64 0.468 ; 
      RECT 3.312 0.252 3.384 0.324 ; 
      RECT 3.096 0.54 3.168 0.612 ; 
      RECT 2.88 0.396 2.952 0.468 ; 
      RECT 2.592 0.54 2.664 0.612 ; 
      RECT 2.432 0.396 2.504 0.468 ; 
      RECT 2.2 0.252 2.272 0.324 ; 
      RECT 2.068 0.54 2.14 0.612 ; 
      RECT 1.692 0.108 1.764 0.18 ; 
      RECT 0.828 0.108 0.9 0.18 ; 
  END 
END SDFLx1_ASAP7_6t_SL 


MACRO SDFLx2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN SDFLx2_ASAP7_6t_SL 0 0 ; 
  SIZE 6.048 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 4.824 0.684 5.304 0.756 ; 
        RECT 5.232 0.108 5.304 0.756 ; 
        RECT 5.128 0.108 5.304 0.184 ; 
        RECT 4.824 0.376 4.896 0.756 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.32 0.396 1.54 0.468 ; 
        RECT 1.32 0.248 1.392 0.468 ; 
        RECT 1.148 0.248 1.392 0.324 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.56 0.684 5.76 0.756 ; 
        RECT 5.688 0.108 5.76 0.756 ; 
        RECT 5.5 0.108 5.76 0.18 ; 
    END 
  END QN 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.396 0.74 0.468 ; 
        RECT 0.128 0.684 0.664 0.756 ; 
        RECT 0.592 0.396 0.664 0.756 ; 
        RECT 0.128 0.108 0.276 0.18 ; 
        RECT 0.128 0.108 0.2 0.756 ; 
    END 
  END SE 
  PIN SI 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.672 0.684 1.936 0.756 ; 
        RECT 1.864 0.396 1.936 0.756 ; 
        RECT 1.672 0.396 1.936 0.468 ; 
    END 
  END SI 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 6.048 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 6.048 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 4.608 0.204 4.68 0.632 ; 
      RECT 4.968 0.54 5.132 0.612 ; 
      RECT 4.968 0.204 5.04 0.612 ; 
      RECT 4.608 0.204 5.04 0.276 ; 
      RECT 3.888 0.684 4.16 0.756 ; 
      RECT 3.888 0.108 3.96 0.756 ; 
      RECT 3.74 0.28 3.96 0.352 ; 
      RECT 3.888 0.108 4.16 0.18 ; 
      RECT 3.4 0.68 3.64 0.752 ; 
      RECT 3.568 0.108 3.64 0.752 ; 
      RECT 3.184 0.108 3.64 0.18 ; 
      RECT 3.312 0.252 3.384 0.492 ; 
      RECT 3.264 0.252 3.424 0.324 ; 
      RECT 3.052 0.54 3.208 0.612 ; 
      RECT 3.096 0.376 3.168 0.612 ; 
      RECT 2.736 0.684 3.16 0.756 ; 
      RECT 2.736 0.188 2.808 0.756 ; 
      RECT 2.664 0.308 2.808 0.38 ; 
      RECT 2.736 0.188 3.06 0.26 ; 
      RECT 2.124 0.684 2.504 0.756 ; 
      RECT 2.432 0.108 2.504 0.756 ; 
      RECT 2.34 0.108 2.504 0.18 ; 
      RECT 2.224 0.252 2.296 0.464 ; 
      RECT 2.148 0.252 2.296 0.324 ; 
      RECT 1.464 0.252 2.004 0.324 ; 
      RECT 1.932 0.108 2.004 0.324 ; 
      RECT 1.464 0.16 1.536 0.324 ; 
      RECT 1.932 0.108 2.196 0.18 ; 
      RECT 2.028 0.54 2.176 0.612 ; 
      RECT 2.028 0.408 2.1 0.612 ; 
      RECT 0.828 0.54 0.9 0.712 ; 
      RECT 0.828 0.54 1.764 0.612 ; 
      RECT 0.344 0.54 0.492 0.612 ; 
      RECT 0.344 0.252 0.42 0.612 ; 
      RECT 0.912 0.396 1.196 0.468 ; 
      RECT 0.912 0.252 0.984 0.468 ; 
      RECT 0.344 0.252 0.984 0.324 ; 
      RECT 5.472 0.352 5.544 0.5 ; 
      RECT 4.464 0.232 4.536 0.632 ; 
      RECT 4.032 0.356 4.104 0.504 ; 
      RECT 3.74 0.452 3.812 0.688 ; 
      RECT 2.88 0.38 2.952 0.576 ; 
      RECT 2.592 0.504 2.664 0.688 ; 
      RECT 1.66 0.108 1.808 0.18 ; 
      RECT 1.044 0.684 1.548 0.756 ; 
      RECT 0.792 0.108 0.94 0.18 ; 
    LAYER M2 ; 
      RECT 3.548 0.396 5.564 0.468 ; 
      RECT 2.048 0.54 4.7 0.612 ; 
      RECT 2.18 0.252 4.556 0.324 ; 
      RECT 2.432 0.396 2.952 0.468 ; 
      RECT 0.768 0.108 1.86 0.18 ; 
    LAYER V1 ; 
      RECT 5.472 0.396 5.544 0.468 ; 
      RECT 4.608 0.54 4.68 0.612 ; 
      RECT 4.464 0.252 4.536 0.324 ; 
      RECT 4.032 0.396 4.104 0.468 ; 
      RECT 3.74 0.54 3.812 0.612 ; 
      RECT 3.568 0.396 3.64 0.468 ; 
      RECT 3.312 0.252 3.384 0.324 ; 
      RECT 3.096 0.54 3.168 0.612 ; 
      RECT 2.88 0.396 2.952 0.468 ; 
      RECT 2.592 0.54 2.664 0.612 ; 
      RECT 2.432 0.396 2.504 0.468 ; 
      RECT 2.2 0.252 2.272 0.324 ; 
      RECT 2.068 0.54 2.14 0.612 ; 
      RECT 1.692 0.108 1.764 0.18 ; 
      RECT 0.828 0.108 0.9 0.18 ; 
  END 
END SDFLx2_ASAP7_6t_SL 


MACRO SDFLx3_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN SDFLx3_ASAP7_6t_SL 0 0 ; 
  SIZE 6.264 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 4.824 0.684 5.304 0.756 ; 
        RECT 5.232 0.108 5.304 0.756 ; 
        RECT 5.128 0.108 5.304 0.184 ; 
        RECT 4.824 0.376 4.896 0.756 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.32 0.396 1.54 0.468 ; 
        RECT 1.32 0.248 1.392 0.468 ; 
        RECT 1.148 0.248 1.392 0.324 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.56 0.684 6.192 0.756 ; 
        RECT 6.12 0.108 6.192 0.756 ; 
        RECT 5.5 0.108 6.192 0.18 ; 
    END 
  END QN 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.396 0.74 0.468 ; 
        RECT 0.128 0.684 0.664 0.756 ; 
        RECT 0.592 0.396 0.664 0.756 ; 
        RECT 0.128 0.108 0.276 0.18 ; 
        RECT 0.128 0.108 0.2 0.756 ; 
    END 
  END SE 
  PIN SI 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.672 0.684 1.936 0.756 ; 
        RECT 1.864 0.396 1.936 0.756 ; 
        RECT 1.672 0.396 1.936 0.468 ; 
    END 
  END SI 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 6.264 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 6.264 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 4.608 0.204 4.68 0.632 ; 
      RECT 4.968 0.54 5.132 0.612 ; 
      RECT 4.968 0.204 5.04 0.612 ; 
      RECT 4.608 0.204 5.04 0.276 ; 
      RECT 3.888 0.684 4.16 0.756 ; 
      RECT 3.888 0.108 3.96 0.756 ; 
      RECT 3.74 0.28 3.96 0.352 ; 
      RECT 3.888 0.108 4.16 0.18 ; 
      RECT 3.4 0.68 3.64 0.752 ; 
      RECT 3.568 0.108 3.64 0.752 ; 
      RECT 3.184 0.108 3.64 0.18 ; 
      RECT 3.312 0.252 3.384 0.492 ; 
      RECT 3.264 0.252 3.424 0.324 ; 
      RECT 3.052 0.54 3.208 0.612 ; 
      RECT 3.096 0.376 3.168 0.612 ; 
      RECT 2.736 0.684 3.16 0.756 ; 
      RECT 2.736 0.188 2.808 0.756 ; 
      RECT 2.664 0.308 2.808 0.38 ; 
      RECT 2.736 0.188 3.06 0.26 ; 
      RECT 2.124 0.684 2.504 0.756 ; 
      RECT 2.432 0.108 2.504 0.756 ; 
      RECT 2.34 0.108 2.504 0.18 ; 
      RECT 2.224 0.252 2.296 0.464 ; 
      RECT 2.148 0.252 2.296 0.324 ; 
      RECT 1.464 0.252 2.004 0.324 ; 
      RECT 1.932 0.108 2.004 0.324 ; 
      RECT 1.464 0.16 1.536 0.324 ; 
      RECT 1.932 0.108 2.196 0.18 ; 
      RECT 2.028 0.54 2.176 0.612 ; 
      RECT 2.028 0.408 2.1 0.612 ; 
      RECT 0.828 0.54 0.9 0.712 ; 
      RECT 0.828 0.54 1.764 0.612 ; 
      RECT 0.344 0.54 0.492 0.612 ; 
      RECT 0.344 0.252 0.42 0.612 ; 
      RECT 0.912 0.396 1.196 0.468 ; 
      RECT 0.912 0.252 0.984 0.468 ; 
      RECT 0.344 0.252 0.984 0.324 ; 
      RECT 5.432 0.396 6.008 0.468 ; 
      RECT 4.464 0.232 4.536 0.632 ; 
      RECT 4.032 0.356 4.104 0.504 ; 
      RECT 3.74 0.452 3.812 0.688 ; 
      RECT 2.88 0.38 2.952 0.576 ; 
      RECT 2.592 0.504 2.664 0.688 ; 
      RECT 1.66 0.108 1.808 0.18 ; 
      RECT 1.044 0.684 1.548 0.756 ; 
      RECT 0.792 0.108 0.94 0.18 ; 
    LAYER M2 ; 
      RECT 3.548 0.396 5.564 0.468 ; 
      RECT 2.048 0.54 4.7 0.612 ; 
      RECT 2.18 0.252 4.556 0.324 ; 
      RECT 2.432 0.396 2.952 0.468 ; 
      RECT 0.768 0.108 1.86 0.18 ; 
    LAYER V1 ; 
      RECT 5.472 0.396 5.544 0.468 ; 
      RECT 4.608 0.54 4.68 0.612 ; 
      RECT 4.464 0.252 4.536 0.324 ; 
      RECT 4.032 0.396 4.104 0.468 ; 
      RECT 3.74 0.54 3.812 0.612 ; 
      RECT 3.568 0.396 3.64 0.468 ; 
      RECT 3.312 0.252 3.384 0.324 ; 
      RECT 3.096 0.54 3.168 0.612 ; 
      RECT 2.88 0.396 2.952 0.468 ; 
      RECT 2.592 0.54 2.664 0.612 ; 
      RECT 2.432 0.396 2.504 0.468 ; 
      RECT 2.2 0.252 2.272 0.324 ; 
      RECT 2.068 0.54 2.14 0.612 ; 
      RECT 1.692 0.108 1.764 0.18 ; 
      RECT 0.828 0.108 0.9 0.18 ; 
  END 
END SDFLx3_ASAP7_6t_SL 


MACRO SDFLx4_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN SDFLx4_ASAP7_6t_SL 0 0 ; 
  SIZE 6.48 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 4.824 0.684 5.304 0.756 ; 
        RECT 5.232 0.108 5.304 0.756 ; 
        RECT 5.128 0.108 5.304 0.184 ; 
        RECT 4.824 0.376 4.896 0.756 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.32 0.396 1.54 0.468 ; 
        RECT 1.32 0.248 1.392 0.468 ; 
        RECT 1.148 0.248 1.392 0.324 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.56 0.684 6.304 0.756 ; 
        RECT 6.232 0.108 6.304 0.756 ; 
        RECT 5.56 0.108 6.304 0.18 ; 
    END 
  END QN 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.396 0.74 0.468 ; 
        RECT 0.128 0.684 0.664 0.756 ; 
        RECT 0.592 0.396 0.664 0.756 ; 
        RECT 0.128 0.108 0.276 0.18 ; 
        RECT 0.128 0.108 0.2 0.756 ; 
    END 
  END SE 
  PIN SI 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.672 0.684 1.936 0.756 ; 
        RECT 1.864 0.396 1.936 0.756 ; 
        RECT 1.672 0.396 1.936 0.468 ; 
    END 
  END SI 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 6.48 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 6.48 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 4.608 0.204 4.68 0.632 ; 
      RECT 4.968 0.54 5.132 0.612 ; 
      RECT 4.968 0.204 5.04 0.612 ; 
      RECT 4.608 0.204 5.04 0.276 ; 
      RECT 3.888 0.684 4.16 0.756 ; 
      RECT 3.888 0.108 3.96 0.756 ; 
      RECT 3.74 0.28 3.96 0.352 ; 
      RECT 3.888 0.108 4.16 0.18 ; 
      RECT 3.4 0.68 3.64 0.752 ; 
      RECT 3.568 0.108 3.64 0.752 ; 
      RECT 3.184 0.108 3.64 0.18 ; 
      RECT 3.312 0.252 3.384 0.492 ; 
      RECT 3.264 0.252 3.424 0.324 ; 
      RECT 3.052 0.54 3.208 0.612 ; 
      RECT 3.096 0.376 3.168 0.612 ; 
      RECT 2.736 0.684 3.16 0.756 ; 
      RECT 2.736 0.188 2.808 0.756 ; 
      RECT 2.664 0.308 2.808 0.38 ; 
      RECT 2.736 0.188 3.06 0.26 ; 
      RECT 2.124 0.684 2.504 0.756 ; 
      RECT 2.432 0.108 2.504 0.756 ; 
      RECT 2.34 0.108 2.504 0.18 ; 
      RECT 2.224 0.252 2.296 0.464 ; 
      RECT 2.148 0.252 2.296 0.324 ; 
      RECT 1.464 0.252 2.004 0.324 ; 
      RECT 1.932 0.108 2.004 0.324 ; 
      RECT 1.464 0.16 1.536 0.324 ; 
      RECT 1.932 0.108 2.196 0.18 ; 
      RECT 2.028 0.54 2.176 0.612 ; 
      RECT 2.028 0.408 2.1 0.612 ; 
      RECT 0.828 0.54 0.9 0.712 ; 
      RECT 0.828 0.54 1.764 0.612 ; 
      RECT 0.344 0.54 0.492 0.612 ; 
      RECT 0.344 0.252 0.42 0.612 ; 
      RECT 0.912 0.396 1.196 0.468 ; 
      RECT 0.912 0.252 0.984 0.468 ; 
      RECT 0.344 0.252 0.984 0.324 ; 
      RECT 5.452 0.396 6.104 0.468 ; 
      RECT 4.464 0.232 4.536 0.632 ; 
      RECT 4.032 0.356 4.104 0.504 ; 
      RECT 3.74 0.452 3.812 0.688 ; 
      RECT 2.88 0.38 2.952 0.576 ; 
      RECT 2.592 0.504 2.664 0.688 ; 
      RECT 1.66 0.108 1.808 0.18 ; 
      RECT 1.044 0.684 1.548 0.756 ; 
      RECT 0.792 0.108 0.94 0.18 ; 
    LAYER M2 ; 
      RECT 3.548 0.396 5.564 0.468 ; 
      RECT 2.048 0.54 4.7 0.612 ; 
      RECT 2.18 0.252 4.556 0.324 ; 
      RECT 2.432 0.396 2.952 0.468 ; 
      RECT 0.768 0.108 1.86 0.18 ; 
    LAYER V1 ; 
      RECT 5.472 0.396 5.544 0.468 ; 
      RECT 4.608 0.54 4.68 0.612 ; 
      RECT 4.464 0.252 4.536 0.324 ; 
      RECT 4.032 0.396 4.104 0.468 ; 
      RECT 3.74 0.54 3.812 0.612 ; 
      RECT 3.568 0.396 3.64 0.468 ; 
      RECT 3.312 0.252 3.384 0.324 ; 
      RECT 3.096 0.54 3.168 0.612 ; 
      RECT 2.88 0.396 2.952 0.468 ; 
      RECT 2.592 0.54 2.664 0.612 ; 
      RECT 2.432 0.396 2.504 0.468 ; 
      RECT 2.2 0.252 2.272 0.324 ; 
      RECT 2.068 0.54 2.14 0.612 ; 
      RECT 1.692 0.108 1.764 0.18 ; 
      RECT 0.828 0.108 0.9 0.18 ; 
  END 
END SDFLx4_ASAP7_6t_SL 


MACRO TAPCELL_ASAP7_6t_SL 
  CLASS CORE WELLTAP ; 
  ORIGIN 0 0 ; 
  FOREIGN TAPCELL_ASAP7_6t_SL 0 0 ; 
  SIZE 0.432 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 0.432 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.432 0.036 ; 
    END 
  END VSS 
END TAPCELL_ASAP7_6t_SL 


MACRO TAPCELL_WITH_FILLER_ASAP7_6t_SL 
  CLASS CORE WELLTAP ; 
  ORIGIN 0 0 ; 
  FOREIGN TAPCELL_WITH_FILLER_ASAP7_6t_SL 0 0 ; 
  SIZE 0.648 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 0.648 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.648 0.036 ; 
    END 
  END VSS 
END TAPCELL_WITH_FILLER_ASAP7_6t_SL 


MACRO TIEHIxp5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN TIEHIxp5_ASAP7_6t_SL 0 0 ; 
  SIZE 0.648 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN H 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.576 0.756 ; 
        RECT 0.504 0.108 0.576 0.756 ; 
        RECT 0.268 0.288 0.576 0.36 ; 
        RECT 0.376 0.108 0.576 0.18 ; 
    END 
  END H 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 0.648 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.648 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 0.072 0.512 0.38 0.584 ; 
      RECT 0.072 0.108 0.144 0.584 ; 
      RECT 0.072 0.108 0.252 0.18 ; 
  END 
END TIEHIxp5_ASAP7_6t_SL 


MACRO TIELOxp5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN TIELOxp5_ASAP7_6t_SL 0 0 ; 
  SIZE 0.648 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN L 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.684 0.576 0.756 ; 
        RECT 0.504 0.108 0.576 0.756 ; 
        RECT 0.268 0.504 0.576 0.576 ; 
        RECT 0.376 0.108 0.576 0.18 ; 
    END 
  END L 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 0.648 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.648 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 0.072 0.684 0.252 0.756 ; 
      RECT 0.072 0.28 0.144 0.756 ; 
      RECT 0.072 0.28 0.38 0.352 ; 
  END 
END TIELOxp5_ASAP7_6t_SL 


MACRO XNOR2x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2x2_ASAP7_6t_SL 0 0 ; 
  SIZE 2.808 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.224 0.396 0.576 0.468 ; 
        RECT 0.32 0.252 0.488 0.468 ; 
        RECT 0.224 0.288 0.38 0.612 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.828 0.396 1.44 0.468 ; 
        RECT 0.072 0.684 0.9 0.756 ; 
        RECT 0.828 0.396 0.9 0.756 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.808 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.808 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.32 0.684 2.52 0.756 ; 
        RECT 2.448 0.108 2.52 0.756 ; 
        RECT 2.26 0.108 2.52 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.692 0.684 1.872 0.756 ; 
      RECT 1.8 0.108 1.872 0.756 ; 
      RECT 1.8 0.4 2.304 0.472 ; 
      RECT 1.392 0.108 1.872 0.18 ; 
      RECT 0.504 0.54 0.756 0.612 ; 
      RECT 0.684 0.108 0.756 0.612 ; 
      RECT 1.584 0.252 1.656 0.488 ; 
      RECT 0.684 0.252 1.656 0.324 ; 
      RECT 0.396 0.108 0.756 0.18 ; 
      RECT 1.024 0.684 1.548 0.756 ; 
  END 
END XNOR2x2_ASAP7_6t_SL 


MACRO XNOR2xp5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2xp5_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.224 0.396 0.576 0.468 ; 
        RECT 0.304 0.396 0.456 0.612 ; 
        RECT 0.224 0.252 0.372 0.468 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.828 0.396 1.44 0.468 ; 
        RECT 0.828 0.108 0.9 0.468 ; 
        RECT 0.072 0.108 0.9 0.18 ; 
        RECT 0.072 0.684 0.22 0.756 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.684 1.872 0.756 ; 
        RECT 1.8 0.108 1.872 0.756 ; 
        RECT 1.692 0.108 1.872 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.684 0.72 0.756 ; 
      RECT 0.648 0.54 0.72 0.756 ; 
      RECT 0.648 0.54 1.656 0.612 ; 
      RECT 1.584 0.376 1.656 0.612 ; 
      RECT 0.684 0.252 0.756 0.612 ; 
      RECT 0.504 0.252 0.756 0.324 ; 
      RECT 1.024 0.108 1.548 0.18 ; 
  END 
END XNOR2xp5_ASAP7_6t_SL 


MACRO XNOR2xp5f_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2xp5f_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.224 0.396 0.576 0.468 ; 
        RECT 0.324 0.396 0.472 0.612 ; 
        RECT 0.224 0.252 0.372 0.468 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.828 0.396 1.44 0.468 ; 
        RECT 0.828 0.108 0.9 0.468 ; 
        RECT 0.072 0.108 0.9 0.18 ; 
        RECT 0.072 0.684 0.272 0.756 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.684 1.872 0.756 ; 
        RECT 1.8 0.108 1.872 0.756 ; 
        RECT 1.672 0.108 1.872 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.396 0.684 0.756 0.756 ; 
      RECT 0.684 0.252 0.756 0.756 ; 
      RECT 0.684 0.54 1.656 0.612 ; 
      RECT 1.584 0.376 1.656 0.612 ; 
      RECT 0.504 0.252 0.756 0.324 ; 
      RECT 1.024 0.108 1.548 0.18 ; 
  END 
END XNOR2xp5f_ASAP7_6t_SL 


MACRO XOR2x2_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2x2_ASAP7_6t_SL 0 0 ; 
  SIZE 2.808 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.224 0.396 0.576 0.468 ; 
        RECT 0.332 0.396 0.48 0.612 ; 
        RECT 0.224 0.252 0.38 0.472 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.828 0.396 1.44 0.468 ; 
        RECT 0.828 0.108 0.9 0.468 ; 
        RECT 0.072 0.108 0.9 0.18 ; 
        RECT 0.072 0.684 0.272 0.756 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 2.808 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.808 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.32 0.684 2.52 0.756 ; 
        RECT 2.448 0.108 2.52 0.756 ; 
        RECT 2.32 0.108 2.52 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.456 0.684 1.872 0.756 ; 
      RECT 1.8 0.108 1.872 0.756 ; 
      RECT 1.8 0.392 2.304 0.464 ; 
      RECT 1.692 0.108 1.872 0.18 ; 
      RECT 0.396 0.684 0.756 0.756 ; 
      RECT 0.684 0.252 0.756 0.756 ; 
      RECT 0.684 0.54 1.656 0.612 ; 
      RECT 1.584 0.376 1.656 0.612 ; 
      RECT 0.504 0.252 0.756 0.324 ; 
      RECT 1.024 0.108 1.568 0.18 ; 
  END 
END XOR2x2_ASAP7_6t_SL 


MACRO XOR2xp5_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2xp5_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.828 0.396 1.44 0.468 ; 
        RECT 0.072 0.684 0.9 0.756 ; 
        RECT 0.828 0.396 0.9 0.756 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.224 0.396 0.576 0.468 ; 
        RECT 0.308 0.252 0.488 0.468 ; 
        RECT 0.224 0.396 0.372 0.612 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.692 0.684 1.872 0.756 ; 
        RECT 1.8 0.108 1.872 0.756 ; 
        RECT 1.024 0.108 1.872 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.504 0.54 0.756 0.612 ; 
      RECT 0.684 0.108 0.756 0.612 ; 
      RECT 1.584 0.252 1.656 0.488 ; 
      RECT 0.684 0.252 1.656 0.324 ; 
      RECT 0.396 0.108 0.756 0.18 ; 
      RECT 1.024 0.684 1.548 0.756 ; 
  END 
END XOR2xp5_ASAP7_6t_SL 


MACRO XOR2xp5r_ASAP7_6t_SL 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2xp5r_ASAP7_6t_SL 0 0 ; 
  SIZE 1.944 BY 0.864 ; 
  SYMMETRY X Y ; 
  SITE asap7sc6t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.224 0.396 0.576 0.468 ; 
        RECT 0.304 0.252 0.456 0.468 ; 
        RECT 0.224 0.396 0.372 0.612 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.828 0.396 1.44 0.468 ; 
        RECT 0.072 0.684 0.9 0.756 ; 
        RECT 0.828 0.396 0.9 0.756 ; 
        RECT 0.072 0.108 0.26 0.18 ; 
        RECT 0.072 0.108 0.144 0.756 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 0.828 1.944 0.9 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.692 0.684 1.872 0.756 ; 
        RECT 1.8 0.108 1.872 0.756 ; 
        RECT 1.024 0.108 1.872 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.504 0.54 0.756 0.612 ; 
      RECT 0.684 0.108 0.756 0.612 ; 
      RECT 1.584 0.252 1.656 0.488 ; 
      RECT 0.684 0.252 1.656 0.324 ; 
      RECT 0.396 0.108 0.756 0.18 ; 
      RECT 1.024 0.684 1.568 0.756 ; 
  END 
END XOR2xp5r_ASAP7_6t_SL 


END LIBRARY 
