# BSD 3-Clause License
# 
# Copyright 2021 Lawrence T. Clark, Vinay Vashishtha, or Arizona State
# University
# 
# Redistribution and use in source and binary forms, with or without
# modification, are permitted provided that the following conditions are met:
# 
# 1. Redistributions of source code must retain the above copyright notice,
# this list of conditions and the following disclaimer.
# 
# 2. Redistributions in binary form must reproduce the above copyright
# notice, this list of conditions and the following disclaimer in the
# documentation and/or other materials provided with the distribution.
# 
# 3. Neither the name of the copyright holder nor the names of its
# contributors may be used to endorse or promote products derived from this
# software without specific prior written permission.
# 
# THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
# AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
# IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
# ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE
# LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
# CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
# SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
# INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
# CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
# ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
# POSSIBILITY OF SUCH DAMAGE.

VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

SITE asap7sc6t
 CLASS CORE ;
 SIZE 0.054 BY 0.216 ;
 SYMMETRY Y ;
END asap7sc6t

MACRO A2O1A1Ixp33_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN A2O1A1Ixp33_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.116 0.056 0.153 ;
        RECT 0.018 0.027 0.036 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1 0.099 0.142 0.117 ;
        RECT 0.081 0.116 0.118 0.153 ;
        RECT 0.1 0.063 0.118 0.153 ;
        RECT 0.081 0.063 0.118 0.081 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.154 0.135 0.195 0.153 ;
        RECT 0.177 0.063 0.195 0.153 ;
        RECT 0.154 0.063 0.195 0.081 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.22 0.135 0.267 0.153 ;
        RECT 0.249 0.08 0.267 0.153 ;
        RECT 0.215 0.063 0.252 0.1 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.171 0.315 0.189 ;
        RECT 0.297 0.027 0.315 0.189 ;
        RECT 0.261 0.027 0.315 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.099 0.027 0.225 0.045 ;
      RECT 0.04 0.171 0.171 0.189 ;
  END
END A2O1A1Ixp33_ASAP7_6t_SL

MACRO A2O1A1Ixp5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN A2O1A1Ixp5_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.135 0.252 0.153 ;
        RECT 0.234 0.106 0.252 0.153 ;
        RECT 0.018 0.171 0.077 0.189 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.067 0.099 0.176 0.117 ;
        RECT 0.067 0.063 0.122 0.081 ;
        RECT 0.067 0.063 0.085 0.117 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.063 0.343 0.081 ;
        RECT 0.288 0.099 0.324 0.117 ;
        RECT 0.306 0.063 0.324 0.117 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.341 0.135 0.378 0.153 ;
        RECT 0.36 0.099 0.378 0.153 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.315 0.171 0.414 0.189 ;
        RECT 0.396 0.027 0.414 0.189 ;
        RECT 0.369 0.027 0.414 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.153 0.063 0.274 0.081 ;
      RECT 0.256 0.027 0.274 0.081 ;
      RECT 0.256 0.027 0.338 0.045 ;
      RECT 0.148 0.171 0.284 0.189 ;
      RECT 0.094 0.027 0.225 0.045 ;
  END
END A2O1A1Ixp5_ASAP7_6t_SL

MACRO A2O1A1O1Ixp33_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN A2O1A1O1Ixp33_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.135 0.055 0.153 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.105 0.099 0.144 0.117 ;
        RECT 0.086 0.134 0.123 0.152 ;
        RECT 0.105 0.063 0.123 0.152 ;
        RECT 0.086 0.063 0.123 0.081 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.135 0.218 0.153 ;
        RECT 0.18 0.063 0.218 0.081 ;
        RECT 0.18 0.063 0.198 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.287 0.135 0.325 0.153 ;
        RECT 0.287 0.063 0.325 0.081 ;
        RECT 0.287 0.063 0.305 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.134 0.414 0.152 ;
        RECT 0.396 0.063 0.414 0.152 ;
        RECT 0.376 0.063 0.414 0.081 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.423 0.171 0.468 0.189 ;
        RECT 0.45 0.027 0.468 0.189 ;
        RECT 0.261 0.027 0.468 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.202 0.171 0.392 0.189 ;
      RECT 0.094 0.027 0.23 0.045 ;
      RECT 0.04 0.171 0.171 0.189 ;
  END
END A2O1A1O1Ixp33_ASAP7_6t_SL

MACRO AND2x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.104 0.135 0.141 0.153 ;
        RECT 0.123 0.063 0.141 0.153 ;
        RECT 0.104 0.063 0.141 0.081 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.09 0.117 ;
        RECT 0.018 0.171 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.171 0.306 0.189 ;
        RECT 0.288 0.027 0.306 0.189 ;
        RECT 0.202 0.027 0.306 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.099 0.171 0.177 0.189 ;
      RECT 0.159 0.027 0.177 0.189 ;
      RECT 0.159 0.099 0.226 0.117 ;
      RECT 0.099 0.027 0.177 0.045 ;
  END
END AND2x2_ASAP7_6t_SL

MACRO AND2x4_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2x4_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.027 0.252 0.117 ;
        RECT 0.018 0.027 0.252 0.045 ;
        RECT 0.018 0.171 0.068 0.189 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.101 0.143 0.119 ;
        RECT 0.088 0.135 0.125 0.153 ;
        RECT 0.107 0.063 0.125 0.153 ;
        RECT 0.088 0.063 0.125 0.081 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.315 0.171 0.522 0.189 ;
        RECT 0.504 0.027 0.522 0.189 ;
        RECT 0.315 0.027 0.522 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.099 0.171 0.283 0.189 ;
      RECT 0.265 0.133 0.283 0.189 ;
      RECT 0.189 0.063 0.207 0.189 ;
      RECT 0.265 0.133 0.306 0.151 ;
      RECT 0.288 0.085 0.306 0.151 ;
      RECT 0.153 0.063 0.207 0.081 ;
  END
END AND2x4_ASAP7_6t_SL

MACRO AND2x6_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2x6_ASAP7_6t_SL 0 0 ;
  SIZE 0.648 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.232 0.027 0.25 0.122 ;
        RECT 0.018 0.027 0.25 0.045 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.135 0.162 0.153 ;
        RECT 0.144 0.099 0.162 0.153 ;
        RECT 0.107 0.099 0.162 0.117 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.648 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.31 0.171 0.63 0.189 ;
        RECT 0.612 0.027 0.63 0.189 ;
        RECT 0.31 0.027 0.63 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.171 0.285 0.189 ;
      RECT 0.267 0.133 0.285 0.189 ;
      RECT 0.18 0.063 0.198 0.189 ;
      RECT 0.267 0.133 0.306 0.151 ;
      RECT 0.288 0.085 0.306 0.151 ;
      RECT 0.115 0.063 0.198 0.081 ;
  END
END AND2x6_ASAP7_6t_SL

MACRO AND3x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.135 0.055 0.153 ;
        RECT 0.018 0.027 0.036 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.099 0.144 0.117 ;
        RECT 0.088 0.135 0.125 0.153 ;
        RECT 0.107 0.027 0.125 0.153 ;
        RECT 0.088 0.027 0.125 0.064 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.161 0.135 0.198 0.153 ;
        RECT 0.18 0.063 0.198 0.153 ;
        RECT 0.161 0.063 0.198 0.081 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.171 0.306 0.189 ;
        RECT 0.288 0.027 0.306 0.189 ;
        RECT 0.261 0.027 0.306 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.171 0.234 0.189 ;
      RECT 0.216 0.027 0.234 0.189 ;
      RECT 0.216 0.099 0.262 0.117 ;
      RECT 0.153 0.027 0.234 0.045 ;
  END
END AND3x1_ASAP7_6t_SL

MACRO AND3x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.135 0.055 0.153 ;
        RECT 0.018 0.027 0.036 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.105 0.099 0.143 0.117 ;
        RECT 0.086 0.135 0.123 0.153 ;
        RECT 0.105 0.027 0.123 0.153 ;
        RECT 0.086 0.027 0.123 0.064 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.158 0.135 0.195 0.153 ;
        RECT 0.177 0.063 0.195 0.153 ;
        RECT 0.158 0.063 0.195 0.081 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.171 0.36 0.189 ;
        RECT 0.342 0.027 0.36 0.189 ;
        RECT 0.256 0.027 0.36 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.171 0.231 0.189 ;
      RECT 0.213 0.027 0.231 0.189 ;
      RECT 0.213 0.099 0.284 0.117 ;
      RECT 0.148 0.027 0.231 0.045 ;
  END
END AND3x2_ASAP7_6t_SL

MACRO AND3x4_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3x4_ASAP7_6t_SL 0 0 ;
  SIZE 0.756 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.688 0.152 0.739 0.189 ;
        RECT 0.721 0.063 0.739 0.189 ;
        RECT 0.702 0.063 0.739 0.081 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.392 0.135 0.567 0.153 ;
        RECT 0.549 0.099 0.567 0.153 ;
        RECT 0.392 0.099 0.567 0.117 ;
        RECT 0.392 0.063 0.429 0.117 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.31 0.135 0.36 0.153 ;
        RECT 0.342 0.081 0.36 0.153 ;
        RECT 0.267 0.081 0.36 0.099 ;
        RECT 0.267 0.027 0.285 0.099 ;
        RECT 0.248 0.027 0.285 0.045 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.756 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.756 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.171 0.212 0.189 ;
        RECT 0.194 0.143 0.212 0.189 ;
        RECT 0.194 0.027 0.212 0.069 ;
        RECT 0.018 0.027 0.212 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.472 0.063 0.603 0.081 ;
      RECT 0.585 0.027 0.603 0.081 ;
      RECT 0.585 0.027 0.718 0.045 ;
      RECT 0.23 0.171 0.646 0.189 ;
      RECT 0.628 0.063 0.646 0.189 ;
      RECT 0.23 0.094 0.248 0.189 ;
      RECT 0.628 0.063 0.67 0.081 ;
      RECT 0.31 0.027 0.554 0.045 ;
  END
END AND3x4_ASAP7_6t_SL

MACRO AND4x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.009 0.152 0.063 0.189 ;
        RECT 0.009 0.028 0.063 0.065 ;
        RECT 0.009 0.099 0.052 0.117 ;
        RECT 0.009 0.028 0.027 0.189 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.081 0.099 0.147 0.117 ;
        RECT 0.081 0.099 0.118 0.153 ;
        RECT 0.081 0.027 0.118 0.064 ;
        RECT 0.081 0.027 0.099 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.16 0.135 0.198 0.153 ;
        RECT 0.18 0.063 0.198 0.153 ;
        RECT 0.136 0.063 0.198 0.081 ;
        RECT 0.136 0.027 0.173 0.081 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.227 0.135 0.264 0.153 ;
        RECT 0.227 0.063 0.264 0.081 ;
        RECT 0.235 0.063 0.253 0.153 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.325 0.171 0.392 0.189 ;
        RECT 0.325 0.027 0.392 0.045 ;
        RECT 0.325 0.027 0.343 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.171 0.307 0.189 ;
      RECT 0.289 0.027 0.307 0.189 ;
      RECT 0.207 0.027 0.307 0.045 ;
  END
END AND4x1_ASAP7_6t_SL

MACRO AND4x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.364 0.171 0.423 0.189 ;
        RECT 0.405 0.028 0.423 0.189 ;
        RECT 0.38 0.099 0.423 0.117 ;
        RECT 0.386 0.028 0.423 0.046 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.318 0.099 0.355 0.153 ;
        RECT 0.337 0.027 0.355 0.153 ;
        RECT 0.311 0.027 0.355 0.064 ;
        RECT 0.283 0.099 0.355 0.117 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.063 0.293 0.081 ;
        RECT 0.256 0.027 0.293 0.081 ;
        RECT 0.234 0.135 0.272 0.153 ;
        RECT 0.234 0.063 0.252 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.166 0.135 0.203 0.153 ;
        RECT 0.166 0.063 0.203 0.081 ;
        RECT 0.179 0.063 0.197 0.153 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.04 0.171 0.105 0.189 ;
        RECT 0.087 0.027 0.105 0.189 ;
        RECT 0.04 0.027 0.105 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.123 0.171 0.333 0.189 ;
      RECT 0.123 0.027 0.141 0.189 ;
      RECT 0.123 0.027 0.225 0.045 ;
  END
END AND4x2_ASAP7_6t_SL

MACRO AND5x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND5x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.027 0.065 0.045 ;
        RECT 0.017 0.027 0.035 0.158 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.103 0.135 0.141 0.153 ;
        RECT 0.123 0.027 0.141 0.153 ;
        RECT 0.097 0.027 0.141 0.045 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.027 0.227 0.045 ;
        RECT 0.159 0.116 0.196 0.153 ;
        RECT 0.178 0.027 0.196 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.252 0.027 0.289 0.052 ;
        RECT 0.231 0.066 0.27 0.084 ;
        RECT 0.252 0.027 0.27 0.084 ;
        RECT 0.214 0.116 0.251 0.153 ;
        RECT 0.231 0.066 0.249 0.153 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.295 0.072 0.339 0.09 ;
        RECT 0.295 0.135 0.334 0.153 ;
        RECT 0.295 0.072 0.313 0.153 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.398 0.027 0.416 0.164 ;
        RECT 0.364 0.027 0.416 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.053 0.171 0.377 0.189 ;
      RECT 0.359 0.096 0.377 0.189 ;
      RECT 0.053 0.091 0.071 0.189 ;
      RECT 0.053 0.091 0.09 0.109 ;
      RECT 0.072 0.066 0.09 0.109 ;
  END
END AND5x1_ASAP7_6t_SL

MACRO AND5x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND5x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.135 0.054 0.153 ;
        RECT 0.036 0.028 0.054 0.153 ;
        RECT 0.017 0.028 0.054 0.046 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.099 0.144 0.117 ;
        RECT 0.072 0.135 0.127 0.153 ;
        RECT 0.072 0.027 0.109 0.045 ;
        RECT 0.072 0.027 0.09 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.063 0.198 0.122 ;
        RECT 0.141 0.027 0.198 0.045 ;
        RECT 0.141 0.063 0.198 0.081 ;
        RECT 0.141 0.027 0.159 0.081 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.135 0.254 0.153 ;
        RECT 0.236 0.081 0.254 0.153 ;
        RECT 0.216 0.063 0.246 0.1 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.282 0.135 0.319 0.153 ;
        RECT 0.282 0.063 0.319 0.081 ;
        RECT 0.288 0.063 0.306 0.153 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.381 0.171 0.468 0.189 ;
        RECT 0.45 0.027 0.468 0.189 ;
        RECT 0.381 0.027 0.468 0.045 ;
        RECT 0.381 0.134 0.399 0.189 ;
        RECT 0.381 0.027 0.399 0.082 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.033 0.171 0.362 0.189 ;
      RECT 0.344 0.027 0.362 0.189 ;
      RECT 0.256 0.027 0.362 0.045 ;
  END
END AND5x2_ASAP7_6t_SL

MACRO AO211x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO211x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.063 0.153 0.081 ;
        RECT 0.129 0.063 0.147 0.12 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.016 0.135 0.053 0.153 ;
        RECT 0.035 0.027 0.053 0.153 ;
        RECT 0.016 0.027 0.053 0.045 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.171 0.284 0.189 ;
        RECT 0.254 0.152 0.284 0.189 ;
        RECT 0.254 0.099 0.272 0.189 ;
        RECT 0.234 0.099 0.272 0.117 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.135 0.223 0.153 ;
        RECT 0.178 0.063 0.216 0.081 ;
        RECT 0.178 0.063 0.196 0.153 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.31 0.171 0.369 0.189 ;
        RECT 0.351 0.027 0.369 0.189 ;
        RECT 0.299 0.027 0.369 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.071 0.135 0.108 0.153 ;
      RECT 0.071 0.027 0.089 0.153 ;
      RECT 0.29 0.063 0.308 0.123 ;
      RECT 0.29 0.099 0.326 0.117 ;
      RECT 0.25 0.063 0.308 0.081 ;
      RECT 0.25 0.027 0.268 0.081 ;
      RECT 0.071 0.027 0.268 0.045 ;
      RECT 0.04 0.171 0.189 0.189 ;
  END
END AO211x1_ASAP7_6t_SL

MACRO AO211x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO211x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.063 0.153 0.081 ;
        RECT 0.129 0.063 0.147 0.132 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.016 0.135 0.053 0.153 ;
        RECT 0.035 0.05 0.053 0.153 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.258 0.14 0.31 0.189 ;
        RECT 0.254 0.099 0.272 0.152 ;
        RECT 0.234 0.099 0.272 0.117 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.063 0.265 0.081 ;
        RECT 0.196 0.171 0.233 0.189 ;
        RECT 0.196 0.134 0.214 0.189 ;
        RECT 0.178 0.063 0.196 0.152 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.328 0.171 0.412 0.189 ;
        RECT 0.394 0.027 0.412 0.189 ;
        RECT 0.328 0.027 0.412 0.045 ;
        RECT 0.328 0.148 0.346 0.189 ;
        RECT 0.328 0.027 0.346 0.069 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.071 0.135 0.108 0.153 ;
      RECT 0.071 0.027 0.089 0.153 ;
      RECT 0.291 0.099 0.346 0.117 ;
      RECT 0.291 0.027 0.309 0.117 ;
      RECT 0.071 0.027 0.309 0.045 ;
      RECT 0.035 0.171 0.171 0.189 ;
  END
END AO211x2_ASAP7_6t_SL

MACRO AO21x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.027 0.068 0.045 ;
        RECT 0.017 0.027 0.035 0.121 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.133 0.135 0.17 0.153 ;
        RECT 0.133 0.063 0.17 0.081 ;
        RECT 0.133 0.063 0.151 0.153 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.201 0.152 0.238 0.189 ;
        RECT 0.201 0.063 0.238 0.1 ;
        RECT 0.201 0.063 0.219 0.189 ;
        RECT 0.183 0.099 0.219 0.117 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.152 0.315 0.189 ;
        RECT 0.297 0.048 0.315 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.071 0.135 0.108 0.153 ;
      RECT 0.071 0.065 0.089 0.153 ;
      RECT 0.261 0.027 0.279 0.122 ;
      RECT 0.071 0.065 0.111 0.083 ;
      RECT 0.093 0.027 0.111 0.083 ;
      RECT 0.093 0.027 0.279 0.045 ;
      RECT 0.04 0.171 0.176 0.189 ;
  END
END AO21x1_ASAP7_6t_SL

MACRO AO21x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.016 0.135 0.053 0.153 ;
        RECT 0.035 0.027 0.053 0.153 ;
        RECT 0.016 0.027 0.053 0.045 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.128 0.063 0.228 0.081 ;
        RECT 0.128 0.135 0.167 0.153 ;
        RECT 0.128 0.063 0.146 0.153 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.182 0.099 0.273 0.117 ;
        RECT 0.207 0.099 0.244 0.189 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.298 0.171 0.362 0.189 ;
        RECT 0.298 0.063 0.323 0.189 ;
        RECT 0.269 0.144 0.323 0.162 ;
        RECT 0.261 0.063 0.323 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.09 0.027 0.108 0.158 ;
      RECT 0.342 0.027 0.36 0.117 ;
      RECT 0.09 0.027 0.36 0.045 ;
      RECT 0.127 0.171 0.182 0.189 ;
      RECT 0.016 0.171 0.068 0.189 ;
    LAYER M2 ;
      RECT 0.04 0.171 0.179 0.189 ;
    LAYER V1 ;
      RECT 0.153 0.171 0.171 0.189 ;
      RECT 0.045 0.171 0.063 0.189 ;
  END
END AO21x2_ASAP7_6t_SL

MACRO AO221x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO221x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.086 0.099 0.141 0.117 ;
        RECT 0.086 0.099 0.123 0.153 ;
        RECT 0.086 0.027 0.123 0.064 ;
        RECT 0.086 0.027 0.104 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.135 0.061 0.153 ;
        RECT 0.018 0.027 0.036 0.153 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.364 0.171 0.401 0.189 ;
        RECT 0.364 0.063 0.401 0.081 ;
        RECT 0.364 0.063 0.382 0.189 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.063 0.265 0.081 ;
        RECT 0.209 0.116 0.246 0.153 ;
        RECT 0.228 0.063 0.246 0.153 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.154 0.135 0.191 0.153 ;
        RECT 0.173 0.063 0.191 0.153 ;
        RECT 0.153 0.063 0.191 0.081 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.472 0.171 0.516 0.189 ;
        RECT 0.498 0.027 0.516 0.189 ;
        RECT 0.472 0.027 0.516 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.271 0.135 0.336 0.153 ;
      RECT 0.318 0.027 0.336 0.153 ;
      RECT 0.429 0.099 0.473 0.117 ;
      RECT 0.429 0.027 0.447 0.117 ;
      RECT 0.148 0.027 0.447 0.045 ;
      RECT 0.207 0.171 0.338 0.189 ;
      RECT 0.04 0.171 0.176 0.189 ;
  END
END AO221x1_ASAP7_6t_SL

MACRO AO221x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO221x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.594 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.086 0.099 0.144 0.117 ;
        RECT 0.086 0.099 0.123 0.153 ;
        RECT 0.086 0.027 0.123 0.064 ;
        RECT 0.086 0.027 0.104 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.135 0.061 0.153 ;
        RECT 0.018 0.027 0.036 0.153 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.364 0.171 0.401 0.189 ;
        RECT 0.364 0.063 0.401 0.081 ;
        RECT 0.364 0.063 0.382 0.189 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.228 0.063 0.265 0.081 ;
        RECT 0.209 0.116 0.246 0.153 ;
        RECT 0.228 0.063 0.246 0.153 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.154 0.135 0.191 0.153 ;
        RECT 0.173 0.063 0.191 0.153 ;
        RECT 0.153 0.063 0.191 0.081 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.594 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.472 0.171 0.516 0.189 ;
        RECT 0.498 0.027 0.516 0.189 ;
        RECT 0.472 0.027 0.516 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.271 0.135 0.336 0.153 ;
      RECT 0.318 0.027 0.336 0.153 ;
      RECT 0.429 0.099 0.473 0.117 ;
      RECT 0.429 0.027 0.447 0.117 ;
      RECT 0.148 0.027 0.447 0.045 ;
      RECT 0.207 0.171 0.338 0.189 ;
      RECT 0.04 0.171 0.176 0.189 ;
  END
END AO221x2_ASAP7_6t_SL

MACRO AO222x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO222x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.594 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.024 0.135 0.069 0.153 ;
        RECT 0.051 0.027 0.069 0.153 ;
        RECT 0.024 0.027 0.069 0.045 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.124 0.135 0.167 0.153 ;
        RECT 0.124 0.063 0.167 0.081 ;
        RECT 0.124 0.063 0.142 0.153 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.283 0.099 0.338 0.117 ;
        RECT 0.32 0.063 0.338 0.117 ;
        RECT 0.283 0.063 0.338 0.081 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.177 0.099 0.253 0.117 ;
        RECT 0.235 0.063 0.253 0.117 ;
        RECT 0.198 0.063 0.253 0.081 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.358 0.099 0.414 0.117 ;
        RECT 0.358 0.063 0.414 0.081 ;
        RECT 0.358 0.063 0.376 0.117 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.44 0.063 0.48 0.1 ;
        RECT 0.411 0.135 0.468 0.153 ;
        RECT 0.45 0.063 0.468 0.153 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.594 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.525 0.171 0.585 0.189 ;
        RECT 0.548 0.152 0.585 0.189 ;
        RECT 0.548 0.027 0.585 0.064 ;
        RECT 0.548 0.027 0.566 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.087 0.027 0.105 0.158 ;
      RECT 0.505 0.027 0.523 0.122 ;
      RECT 0.087 0.027 0.523 0.045 ;
      RECT 0.342 0.171 0.468 0.189 ;
      RECT 0.342 0.135 0.36 0.189 ;
      RECT 0.211 0.135 0.36 0.153 ;
      RECT 0.256 0.171 0.309 0.189 ;
      RECT 0.148 0.171 0.185 0.189 ;
      RECT 0.018 0.171 0.068 0.189 ;
    LAYER M2 ;
      RECT 0.02 0.171 0.287 0.189 ;
    LAYER V1 ;
      RECT 0.261 0.171 0.279 0.189 ;
      RECT 0.153 0.171 0.171 0.189 ;
      RECT 0.045 0.171 0.063 0.189 ;
  END
END AO222x1_ASAP7_6t_SL

MACRO AO222x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO222x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.648 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.052 0.099 0.07 0.14 ;
        RECT 0.016 0.027 0.068 0.064 ;
        RECT 0.016 0.099 0.07 0.117 ;
        RECT 0.016 0.027 0.034 0.117 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.124 0.063 0.167 0.081 ;
        RECT 0.124 0.135 0.162 0.153 ;
        RECT 0.124 0.063 0.142 0.153 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.283 0.099 0.338 0.117 ;
        RECT 0.32 0.063 0.338 0.117 ;
        RECT 0.283 0.063 0.338 0.081 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.182 0.099 0.253 0.117 ;
        RECT 0.2 0.065 0.253 0.117 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.358 0.099 0.414 0.117 ;
        RECT 0.358 0.063 0.414 0.081 ;
        RECT 0.358 0.063 0.376 0.117 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.44 0.063 0.482 0.1 ;
        RECT 0.411 0.135 0.468 0.153 ;
        RECT 0.45 0.063 0.468 0.153 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.648 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.526 0.171 0.63 0.189 ;
        RECT 0.612 0.027 0.63 0.189 ;
        RECT 0.544 0.027 0.63 0.045 ;
        RECT 0.544 0.027 0.562 0.074 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.088 0.027 0.106 0.17 ;
      RECT 0.508 0.027 0.526 0.117 ;
      RECT 0.088 0.027 0.526 0.045 ;
      RECT 0.342 0.171 0.468 0.189 ;
      RECT 0.342 0.135 0.36 0.189 ;
      RECT 0.211 0.135 0.36 0.153 ;
      RECT 0.018 0.171 0.065 0.189 ;
      RECT 0.018 0.152 0.036 0.189 ;
      RECT 0.256 0.171 0.309 0.189 ;
      RECT 0.148 0.171 0.185 0.189 ;
    LAYER M2 ;
      RECT 0.02 0.171 0.287 0.189 ;
    LAYER V1 ;
      RECT 0.261 0.171 0.279 0.189 ;
      RECT 0.153 0.171 0.171 0.189 ;
      RECT 0.045 0.171 0.063 0.189 ;
  END
END AO222x2_ASAP7_6t_SL

MACRO AO22x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.031 0.135 0.068 0.153 ;
        RECT 0.05 0.027 0.068 0.153 ;
        RECT 0.031 0.027 0.068 0.045 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.105 0.098 0.141 0.116 ;
        RECT 0.086 0.116 0.123 0.153 ;
        RECT 0.105 0.027 0.123 0.153 ;
        RECT 0.086 0.027 0.123 0.064 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.309 0.171 0.346 0.189 ;
        RECT 0.309 0.063 0.346 0.081 ;
        RECT 0.309 0.063 0.327 0.189 ;
        RECT 0.286 0.099 0.327 0.117 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.155 0.135 0.192 0.153 ;
        RECT 0.174 0.027 0.192 0.153 ;
        RECT 0.148 0.027 0.192 0.065 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.418 0.171 0.458 0.189 ;
        RECT 0.44 0.027 0.458 0.189 ;
        RECT 0.418 0.027 0.458 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.217 0.135 0.254 0.153 ;
      RECT 0.235 0.027 0.254 0.153 ;
      RECT 0.374 0.099 0.415 0.117 ;
      RECT 0.374 0.027 0.392 0.117 ;
      RECT 0.217 0.054 0.254 0.072 ;
      RECT 0.235 0.027 0.392 0.045 ;
      RECT 0.04 0.171 0.284 0.189 ;
  END
END AO22x1_ASAP7_6t_SL

MACRO AO22x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.031 0.135 0.068 0.153 ;
        RECT 0.05 0.027 0.068 0.153 ;
        RECT 0.031 0.027 0.068 0.045 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.105 0.098 0.141 0.116 ;
        RECT 0.086 0.116 0.123 0.153 ;
        RECT 0.105 0.027 0.123 0.153 ;
        RECT 0.086 0.027 0.123 0.064 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.309 0.171 0.346 0.189 ;
        RECT 0.309 0.063 0.346 0.081 ;
        RECT 0.309 0.063 0.327 0.189 ;
        RECT 0.286 0.099 0.327 0.117 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.155 0.135 0.192 0.153 ;
        RECT 0.174 0.027 0.192 0.153 ;
        RECT 0.148 0.027 0.192 0.065 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.418 0.171 0.459 0.189 ;
        RECT 0.441 0.027 0.459 0.189 ;
        RECT 0.418 0.027 0.459 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.217 0.135 0.254 0.153 ;
      RECT 0.235 0.027 0.254 0.153 ;
      RECT 0.374 0.099 0.415 0.117 ;
      RECT 0.374 0.027 0.392 0.117 ;
      RECT 0.217 0.054 0.254 0.072 ;
      RECT 0.235 0.027 0.392 0.045 ;
      RECT 0.04 0.171 0.284 0.189 ;
  END
END AO22x2_ASAP7_6t_SL

MACRO AO311x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO311x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.063 0.222 0.081 ;
        RECT 0.178 0.063 0.196 0.122 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.135 0.144 0.153 ;
        RECT 0.126 0.027 0.144 0.153 ;
        RECT 0.094 0.027 0.144 0.045 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.093 0.117 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.217 0.135 0.254 0.153 ;
        RECT 0.236 0.096 0.254 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.063 0.306 0.146 ;
        RECT 0.269 0.063 0.306 0.081 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.472 0.171 0.521 0.189 ;
        RECT 0.503 0.027 0.521 0.189 ;
        RECT 0.472 0.027 0.521 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.31 0.171 0.36 0.189 ;
      RECT 0.342 0.027 0.36 0.189 ;
      RECT 0.342 0.099 0.471 0.117 ;
      RECT 0.198 0.027 0.36 0.045 ;
      RECT 0.094 0.171 0.234 0.189 ;
  END
END AO311x1_ASAP7_6t_SL

MACRO AO311x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO311x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.594 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.063 0.217 0.081 ;
        RECT 0.18 0.063 0.198 0.122 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.135 0.144 0.153 ;
        RECT 0.126 0.027 0.144 0.153 ;
        RECT 0.094 0.027 0.144 0.045 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.093 0.117 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.217 0.135 0.254 0.153 ;
        RECT 0.236 0.094 0.254 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.29 0.063 0.308 0.146 ;
        RECT 0.271 0.063 0.308 0.081 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.594 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.472 0.171 0.575 0.189 ;
        RECT 0.557 0.027 0.575 0.189 ;
        RECT 0.472 0.027 0.575 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.31 0.171 0.36 0.189 ;
      RECT 0.342 0.027 0.36 0.189 ;
      RECT 0.342 0.099 0.473 0.117 ;
      RECT 0.198 0.027 0.36 0.045 ;
      RECT 0.094 0.171 0.234 0.189 ;
  END
END AO311x2_ASAP7_6t_SL

MACRO AO31x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO31x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.115 0.063 0.153 0.1 ;
        RECT 0.098 0.135 0.141 0.153 ;
        RECT 0.123 0.063 0.141 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.063 0.222 0.081 ;
        RECT 0.174 0.135 0.211 0.153 ;
        RECT 0.178 0.063 0.196 0.153 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.255 0.152 0.292 0.189 ;
        RECT 0.255 0.099 0.273 0.189 ;
        RECT 0.231 0.099 0.273 0.117 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.027 0.054 0.045 ;
        RECT 0.017 0.027 0.035 0.158 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.323 0.171 0.36 0.189 ;
        RECT 0.342 0.027 0.36 0.189 ;
        RECT 0.305 0.027 0.36 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.055 0.074 0.073 0.158 ;
      RECT 0.306 0.063 0.324 0.122 ;
      RECT 0.055 0.074 0.097 0.092 ;
      RECT 0.079 0.027 0.097 0.092 ;
      RECT 0.256 0.063 0.324 0.081 ;
      RECT 0.256 0.027 0.274 0.081 ;
      RECT 0.079 0.027 0.274 0.045 ;
      RECT 0.094 0.171 0.23 0.189 ;
  END
END AO31x1_ASAP7_6t_SL

MACRO AO31x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO31x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.115 0.063 0.152 0.1 ;
        RECT 0.098 0.135 0.141 0.153 ;
        RECT 0.123 0.063 0.141 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.063 0.215 0.081 ;
        RECT 0.166 0.135 0.207 0.153 ;
        RECT 0.178 0.063 0.196 0.153 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.254 0.152 0.31 0.189 ;
        RECT 0.254 0.099 0.272 0.189 ;
        RECT 0.231 0.099 0.272 0.117 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.027 0.054 0.045 ;
        RECT 0.017 0.027 0.035 0.158 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.328 0.171 0.412 0.189 ;
        RECT 0.394 0.027 0.412 0.189 ;
        RECT 0.328 0.027 0.412 0.045 ;
        RECT 0.328 0.148 0.346 0.189 ;
        RECT 0.328 0.027 0.346 0.069 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.055 0.074 0.073 0.158 ;
      RECT 0.29 0.099 0.345 0.117 ;
      RECT 0.29 0.027 0.308 0.117 ;
      RECT 0.055 0.074 0.097 0.092 ;
      RECT 0.079 0.027 0.097 0.092 ;
      RECT 0.079 0.027 0.308 0.045 ;
      RECT 0.094 0.171 0.225 0.189 ;
  END
END AO31x2_ASAP7_6t_SL

MACRO AO321x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO321x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.594 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.594 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.526 0.171 0.575 0.189 ;
        RECT 0.557 0.027 0.575 0.189 ;
        RECT 0.526 0.027 0.575 0.045 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.15 0.099 0.228 0.117 ;
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.122 ;
      LAYER V1 ;
        RECT 0.18 0.099 0.198 0.117 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.091 0.063 0.174 0.081 ;
      LAYER M1 ;
        RECT 0.098 0.135 0.144 0.153 ;
        RECT 0.126 0.027 0.144 0.153 ;
        RECT 0.094 0.027 0.144 0.045 ;
      LAYER V1 ;
        RECT 0.126 0.063 0.144 0.081 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.258 0.063 0.336 0.081 ;
      LAYER M1 ;
        RECT 0.288 0.057 0.306 0.117 ;
      LAYER V1 ;
        RECT 0.288 0.063 0.306 0.081 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.312 0.099 0.39 0.117 ;
      LAYER M1 ;
        RECT 0.339 0.099 0.394 0.117 ;
        RECT 0.339 0.063 0.394 0.081 ;
        RECT 0.339 0.063 0.357 0.117 ;
      LAYER V1 ;
        RECT 0.342 0.099 0.36 0.117 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.204 0.135 0.282 0.153 ;
      LAYER M1 ;
        RECT 0.222 0.135 0.271 0.153 ;
        RECT 0.234 0.07 0.252 0.153 ;
      LAYER V1 ;
        RECT 0.234 0.135 0.252 0.153 ;
    END
  END C
  OBS
    LAYER M1 ;
      RECT 0.315 0.135 0.446 0.153 ;
      RECT 0.428 0.027 0.446 0.153 ;
      RECT 0.428 0.099 0.525 0.117 ;
      RECT 0.35 0.027 0.446 0.045 ;
      RECT 0.261 0.171 0.396 0.189 ;
      RECT 0.198 0.027 0.238 0.045 ;
      RECT 0.094 0.171 0.23 0.189 ;
    LAYER M2 ;
      RECT 0.202 0.027 0.446 0.045 ;
    LAYER V1 ;
      RECT 0.423 0.027 0.441 0.045 ;
      RECT 0.207 0.027 0.225 0.045 ;
  END
END AO321x1_ASAP7_6t_SL

MACRO AO321x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO321x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.648 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.648 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.122 ;
      LAYER M2 ;
        RECT 0.15 0.099 0.228 0.117 ;
      LAYER V1 ;
        RECT 0.18 0.099 0.198 0.117 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.135 0.144 0.153 ;
        RECT 0.126 0.027 0.144 0.153 ;
        RECT 0.094 0.027 0.144 0.045 ;
      LAYER M2 ;
        RECT 0.096 0.063 0.174 0.081 ;
      LAYER V1 ;
        RECT 0.126 0.063 0.144 0.081 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
      LAYER M2 ;
        RECT 0.018 0.135 0.096 0.153 ;
      LAYER V1 ;
        RECT 0.018 0.135 0.036 0.153 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.277 0.027 0.317 0.045 ;
        RECT 0.288 0.027 0.306 0.117 ;
      LAYER M2 ;
        RECT 0.258 0.063 0.336 0.081 ;
      LAYER V1 ;
        RECT 0.288 0.063 0.306 0.081 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.339 0.099 0.397 0.117 ;
        RECT 0.339 0.063 0.397 0.081 ;
        RECT 0.339 0.063 0.357 0.117 ;
      LAYER M2 ;
        RECT 0.33 0.099 0.408 0.117 ;
      LAYER V1 ;
        RECT 0.36 0.099 0.378 0.117 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.135 0.271 0.153 ;
        RECT 0.234 0.07 0.252 0.153 ;
      LAYER M2 ;
        RECT 0.206 0.135 0.284 0.153 ;
      LAYER V1 ;
        RECT 0.236 0.135 0.254 0.153 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.526 0.171 0.629 0.189 ;
        RECT 0.611 0.027 0.629 0.189 ;
        RECT 0.526 0.027 0.629 0.045 ;
      LAYER M2 ;
        RECT 0.551 0.099 0.629 0.117 ;
      LAYER V1 ;
        RECT 0.611 0.099 0.629 0.117 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.315 0.135 0.446 0.153 ;
      RECT 0.428 0.027 0.446 0.153 ;
      RECT 0.428 0.099 0.525 0.117 ;
      RECT 0.356 0.027 0.446 0.045 ;
      RECT 0.256 0.171 0.396 0.189 ;
      RECT 0.198 0.027 0.238 0.045 ;
      RECT 0.094 0.171 0.225 0.189 ;
    LAYER M2 ;
      RECT 0.207 0.027 0.441 0.045 ;
    LAYER V1 ;
      RECT 0.423 0.027 0.441 0.045 ;
      RECT 0.207 0.027 0.225 0.045 ;
  END
END AO321x2_ASAP7_6t_SL

MACRO AO322x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO322x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.648 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.522 0.116 0.559 0.153 ;
        RECT 0.504 0.099 0.555 0.117 ;
        RECT 0.537 0.027 0.555 0.153 ;
        RECT 0.522 0.096 0.555 0.153 ;
        RECT 0.518 0.027 0.555 0.064 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.027 0.5 0.064 ;
        RECT 0.45 0.135 0.487 0.153 ;
        RECT 0.45 0.027 0.468 0.153 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.359 0.135 0.425 0.153 ;
        RECT 0.396 0.027 0.414 0.153 ;
        RECT 0.371 0.027 0.414 0.064 ;
        RECT 0.364 0.027 0.414 0.061 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.209 0.099 0.267 0.117 ;
        RECT 0.249 0.063 0.267 0.117 ;
        RECT 0.208 0.063 0.267 0.081 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.099 0.361 0.117 ;
        RECT 0.285 0.063 0.34 0.081 ;
        RECT 0.285 0.063 0.303 0.117 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.027 0.068 0.064 ;
        RECT 0.009 0.116 0.046 0.153 ;
        RECT 0.017 0.027 0.035 0.153 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.122 0.099 0.178 0.117 ;
        RECT 0.122 0.063 0.177 0.081 ;
        RECT 0.122 0.063 0.14 0.117 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.648 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.613 0.027 0.631 0.179 ;
        RECT 0.58 0.027 0.631 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.526 0.171 0.595 0.189 ;
      RECT 0.577 0.094 0.595 0.189 ;
      RECT 0.032 0.171 0.091 0.189 ;
      RECT 0.072 0.097 0.091 0.189 ;
      RECT 0.086 0.027 0.104 0.115 ;
      RECT 0.086 0.027 0.333 0.045 ;
      RECT 0.109 0.135 0.127 0.176 ;
      RECT 0.109 0.135 0.328 0.153 ;
      RECT 0.261 0.171 0.495 0.189 ;
      RECT 0.193 0.171 0.23 0.189 ;
    LAYER M2 ;
      RECT 0.04 0.171 0.554 0.189 ;
    LAYER V1 ;
      RECT 0.531 0.171 0.549 0.189 ;
      RECT 0.207 0.171 0.225 0.189 ;
      RECT 0.045 0.171 0.063 0.189 ;
  END
END AO322x1_ASAP7_6t_SL

MACRO AO322x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO322x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.702 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.538 0.027 0.617 0.045 ;
        RECT 0.538 0.135 0.579 0.153 ;
        RECT 0.538 0.027 0.556 0.153 ;
        RECT 0.499 0.099 0.556 0.117 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.135 0.505 0.153 ;
        RECT 0.45 0.063 0.505 0.081 ;
        RECT 0.45 0.063 0.468 0.153 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.414 0.027 0.506 0.045 ;
        RECT 0.414 0.027 0.432 0.094 ;
        RECT 0.359 0.135 0.425 0.153 ;
        RECT 0.396 0.067 0.414 0.153 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.214 0.099 0.269 0.117 ;
        RECT 0.251 0.063 0.269 0.117 ;
        RECT 0.214 0.063 0.269 0.081 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.287 0.099 0.361 0.117 ;
        RECT 0.287 0.063 0.342 0.081 ;
        RECT 0.287 0.063 0.305 0.117 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.135 0.054 0.153 ;
        RECT 0.036 0.027 0.054 0.153 ;
        RECT 0.017 0.027 0.054 0.081 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.109 0.099 0.181 0.117 ;
        RECT 0.109 0.063 0.181 0.081 ;
        RECT 0.109 0.063 0.127 0.117 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.702 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.702 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.581 0.063 0.685 0.081 ;
        RECT 0.648 0.027 0.685 0.081 ;
        RECT 0.567 0.171 0.622 0.189 ;
        RECT 0.604 0.063 0.622 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.651 0.171 0.688 0.189 ;
      RECT 0.67 0.099 0.688 0.189 ;
      RECT 0.647 0.099 0.688 0.117 ;
      RECT 0.036 0.171 0.091 0.189 ;
      RECT 0.073 0.027 0.091 0.189 ;
      RECT 0.073 0.027 0.387 0.045 ;
      RECT 0.112 0.135 0.13 0.176 ;
      RECT 0.112 0.135 0.328 0.153 ;
      RECT 0.261 0.171 0.5 0.189 ;
      RECT 0.166 0.171 0.23 0.189 ;
    LAYER M2 ;
      RECT 0.036 0.171 0.682 0.189 ;
    LAYER V1 ;
      RECT 0.657 0.171 0.675 0.189 ;
      RECT 0.207 0.171 0.225 0.189 ;
      RECT 0.045 0.171 0.063 0.189 ;
  END
END AO322x2_ASAP7_6t_SL

MACRO AO32x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO32x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.214 0.116 0.251 0.153 ;
        RECT 0.233 0.027 0.251 0.153 ;
        RECT 0.214 0.027 0.251 0.064 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.159 0.116 0.196 0.153 ;
        RECT 0.178 0.027 0.196 0.153 ;
        RECT 0.153 0.027 0.196 0.045 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.063 0.144 0.081 ;
        RECT 0.123 0.063 0.141 0.153 ;
        RECT 0.099 0.135 0.141 0.153 ;
        RECT 0.085 0.152 0.122 0.189 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.269 0.116 0.306 0.153 ;
        RECT 0.288 0.087 0.306 0.153 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.386 0.027 0.423 0.084 ;
        RECT 0.379 0.135 0.416 0.153 ;
        RECT 0.379 0.064 0.397 0.153 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.023 0.171 0.06 0.189 ;
        RECT 0.023 0.041 0.041 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.324 0.027 0.342 0.16 ;
      RECT 0.301 0.027 0.361 0.045 ;
      RECT 0.064 0.027 0.082 0.117 ;
      RECT 0.064 0.027 0.122 0.045 ;
      RECT 0.363 0.171 0.416 0.189 ;
      RECT 0.153 0.171 0.287 0.189 ;
    LAYER M2 ;
      RECT 0.202 0.171 0.395 0.189 ;
      RECT 0.094 0.027 0.353 0.045 ;
    LAYER V1 ;
      RECT 0.369 0.171 0.387 0.189 ;
      RECT 0.315 0.027 0.333 0.045 ;
      RECT 0.207 0.171 0.225 0.189 ;
      RECT 0.099 0.027 0.117 0.045 ;
  END
END AO32x1_ASAP7_6t_SL

MACRO AO32x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO32x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.268 0.116 0.305 0.153 ;
        RECT 0.287 0.042 0.305 0.153 ;
        RECT 0.268 0.042 0.305 0.079 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.213 0.116 0.25 0.153 ;
        RECT 0.232 0.044 0.25 0.153 ;
        RECT 0.213 0.044 0.25 0.081 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.138 0.135 0.195 0.153 ;
        RECT 0.177 0.058 0.195 0.153 ;
        RECT 0.095 0.171 0.174 0.189 ;
        RECT 0.138 0.135 0.174 0.189 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.323 0.116 0.36 0.153 ;
        RECT 0.342 0.042 0.36 0.153 ;
        RECT 0.323 0.042 0.36 0.079 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.414 0.116 0.47 0.153 ;
        RECT 0.452 0.063 0.47 0.153 ;
        RECT 0.421 0.063 0.47 0.085 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.063 0.112 0.081 ;
        RECT 0.018 0.135 0.107 0.153 ;
        RECT 0.018 0.135 0.055 0.189 ;
        RECT 0.018 0.027 0.055 0.081 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.378 0.027 0.396 0.16 ;
      RECT 0.378 0.027 0.446 0.045 ;
      RECT 0.084 0.099 0.155 0.117 ;
      RECT 0.137 0.027 0.155 0.117 ;
      RECT 0.094 0.027 0.156 0.045 ;
      RECT 0.418 0.171 0.47 0.189 ;
      RECT 0.207 0.171 0.341 0.189 ;
    LAYER M2 ;
      RECT 0.31 0.171 0.449 0.189 ;
      RECT 0.094 0.027 0.446 0.045 ;
    LAYER V1 ;
      RECT 0.423 0.027 0.441 0.045 ;
      RECT 0.423 0.171 0.441 0.189 ;
      RECT 0.315 0.171 0.333 0.189 ;
      RECT 0.099 0.027 0.117 0.045 ;
  END
END AO32x2_ASAP7_6t_SL

MACRO AO331x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO331x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.135 0.271 0.153 ;
        RECT 0.224 0.027 0.261 0.045 ;
        RECT 0.234 0.027 0.252 0.153 ;
      LAYER M2 ;
        RECT 0.205 0.135 0.301 0.153 ;
      LAYER V1 ;
        RECT 0.247 0.135 0.265 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.135 0.208 0.153 ;
        RECT 0.181 0.027 0.199 0.153 ;
        RECT 0.162 0.027 0.199 0.045 ;
      LAYER M2 ;
        RECT 0.131 0.099 0.247 0.117 ;
      LAYER V1 ;
        RECT 0.181 0.099 0.199 0.117 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.104 0.135 0.144 0.153 ;
        RECT 0.126 0.099 0.144 0.153 ;
      LAYER M2 ;
        RECT 0.076 0.135 0.173 0.153 ;
      LAYER V1 ;
        RECT 0.117 0.135 0.135 0.153 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.286 0.027 0.323 0.045 ;
        RECT 0.286 0.027 0.304 0.11 ;
      LAYER M2 ;
        RECT 0.239 0.063 0.355 0.081 ;
      LAYER V1 ;
        RECT 0.286 0.063 0.304 0.081 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.334 0.099 0.371 0.117 ;
        RECT 0.343 0.07 0.361 0.117 ;
      LAYER M2 ;
        RECT 0.293 0.099 0.412 0.117 ;
      LAYER V1 ;
        RECT 0.347 0.099 0.365 0.117 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.063 0.443 0.081 ;
        RECT 0.396 0.063 0.414 0.11 ;
      LAYER M2 ;
        RECT 0.402 0.063 0.511 0.081 ;
      LAYER V1 ;
        RECT 0.423 0.063 0.441 0.081 ;
    END
  END B3
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.452 0.099 0.495 0.117 ;
        RECT 0.477 0.07 0.495 0.117 ;
      LAYER M2 ;
        RECT 0.446 0.099 0.511 0.117 ;
      LAYER V1 ;
        RECT 0.469 0.099 0.487 0.117 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.171 0.068 0.189 ;
        RECT 0.018 0.027 0.063 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
      LAYER M2 ;
        RECT 0.039 0.171 0.137 0.189 ;
      LAYER V1 ;
        RECT 0.045 0.171 0.063 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.452 0.171 0.531 0.189 ;
      RECT 0.513 0.027 0.531 0.189 ;
      RECT 0.364 0.027 0.531 0.045 ;
      RECT 0.072 0.063 0.09 0.117 ;
      RECT 0.072 0.063 0.112 0.081 ;
      RECT 0.094 0.027 0.112 0.081 ;
      RECT 0.094 0.027 0.131 0.045 ;
      RECT 0.315 0.135 0.465 0.153 ;
      RECT 0.138 0.171 0.393 0.189 ;
    LAYER M2 ;
      RECT 0.094 0.027 0.446 0.045 ;
    LAYER V1 ;
      RECT 0.423 0.027 0.441 0.045 ;
      RECT 0.099 0.027 0.117 0.045 ;
  END
END AO331x1_ASAP7_6t_SL

MACRO AO331x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO331x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.594 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.594 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.135 0.327 0.153 ;
        RECT 0.288 0.053 0.306 0.153 ;
      LAYER M2 ;
        RECT 0.263 0.135 0.38 0.153 ;
      LAYER V1 ;
        RECT 0.297 0.135 0.315 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.225 0.135 0.262 0.153 ;
        RECT 0.233 0.053 0.251 0.153 ;
      LAYER M2 ;
        RECT 0.206 0.063 0.28 0.081 ;
      LAYER V1 ;
        RECT 0.233 0.063 0.251 0.081 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.161 0.135 0.198 0.153 ;
        RECT 0.18 0.099 0.198 0.153 ;
      LAYER M2 ;
        RECT 0.113 0.135 0.224 0.153 ;
      LAYER V1 ;
        RECT 0.167 0.135 0.185 0.153 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.336 0.099 0.364 0.117 ;
        RECT 0.34 0.053 0.358 0.117 ;
      LAYER M2 ;
        RECT 0.335 0.099 0.412 0.117 ;
      LAYER V1 ;
        RECT 0.342 0.099 0.36 0.117 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.383 0.063 0.425 0.081 ;
        RECT 0.397 0.063 0.415 0.11 ;
      LAYER M2 ;
        RECT 0.383 0.063 0.453 0.081 ;
      LAYER V1 ;
        RECT 0.388 0.063 0.406 0.081 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.063 0.534 0.081 ;
        RECT 0.45 0.063 0.468 0.11 ;
      LAYER M2 ;
        RECT 0.484 0.063 0.572 0.081 ;
      LAYER V1 ;
        RECT 0.504 0.063 0.522 0.081 ;
    END
  END B3
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.499 0.099 0.542 0.117 ;
      LAYER M2 ;
        RECT 0.484 0.099 0.572 0.117 ;
      LAYER V1 ;
        RECT 0.504 0.099 0.522 0.117 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.171 0.122 0.189 ;
        RECT 0.018 0.027 0.117 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
      LAYER M2 ;
        RECT 0.093 0.171 0.191 0.189 ;
      LAYER V1 ;
        RECT 0.099 0.171 0.117 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.526 0.171 0.585 0.189 ;
      RECT 0.567 0.027 0.585 0.189 ;
      RECT 0.418 0.027 0.585 0.045 ;
      RECT 0.105 0.063 0.123 0.122 ;
      RECT 0.105 0.063 0.168 0.081 ;
      RECT 0.148 0.027 0.168 0.081 ;
      RECT 0.148 0.027 0.185 0.045 ;
      RECT 0.374 0.135 0.5 0.153 ;
      RECT 0.197 0.171 0.447 0.189 ;
    LAYER M2 ;
      RECT 0.148 0.027 0.446 0.045 ;
    LAYER V1 ;
      RECT 0.423 0.027 0.441 0.045 ;
      RECT 0.153 0.027 0.171 0.045 ;
  END
END AO331x2_ASAP7_6t_SL

MACRO AO332x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO332x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.756 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.159 0.097 0.2 0.115 ;
        RECT 0.159 0.027 0.177 0.158 ;
        RECT 0.094 0.027 0.177 0.045 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.135 0.141 0.153 ;
        RECT 0.123 0.063 0.141 0.153 ;
        RECT 0.068 0.063 0.141 0.081 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.212 0.135 0.249 0.153 ;
        RECT 0.231 0.027 0.249 0.153 ;
        RECT 0.202 0.027 0.249 0.045 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.267 0.027 0.338 0.045 ;
        RECT 0.267 0.099 0.322 0.117 ;
        RECT 0.267 0.027 0.285 0.117 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.357 0.099 0.412 0.117 ;
        RECT 0.31 0.063 0.412 0.081 ;
        RECT 0.357 0.063 0.375 0.117 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.171 0.632 0.189 ;
        RECT 0.614 0.063 0.632 0.189 ;
        RECT 0.592 0.063 0.632 0.081 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.445 0.099 0.53 0.117 ;
        RECT 0.512 0.063 0.53 0.117 ;
        RECT 0.445 0.063 0.53 0.081 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.756 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.756 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.688 0.171 0.738 0.189 ;
        RECT 0.72 0.027 0.738 0.189 ;
        RECT 0.701 0.027 0.738 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.482 0.135 0.567 0.153 ;
      RECT 0.549 0.027 0.567 0.153 ;
      RECT 0.65 0.099 0.695 0.117 ;
      RECT 0.65 0.027 0.668 0.117 ;
      RECT 0.369 0.027 0.668 0.045 ;
      RECT 0.433 0.171 0.549 0.189 ;
      RECT 0.433 0.135 0.451 0.189 ;
      RECT 0.275 0.135 0.451 0.153 ;
      RECT 0.193 0.171 0.392 0.189 ;
      RECT 0.094 0.171 0.135 0.189 ;
    LAYER M2 ;
      RECT 0.099 0.171 0.234 0.189 ;
    LAYER V1 ;
      RECT 0.207 0.171 0.225 0.189 ;
      RECT 0.099 0.171 0.117 0.189 ;
  END
END AO332x1_ASAP7_6t_SL

MACRO AO332x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO332x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.81 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.159 0.097 0.2 0.115 ;
        RECT 0.159 0.027 0.177 0.158 ;
        RECT 0.094 0.027 0.177 0.045 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.135 0.141 0.153 ;
        RECT 0.123 0.063 0.141 0.153 ;
        RECT 0.068 0.063 0.141 0.081 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.135 0.249 0.153 ;
        RECT 0.231 0.027 0.249 0.153 ;
        RECT 0.202 0.027 0.249 0.045 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.267 0.027 0.338 0.045 ;
        RECT 0.267 0.099 0.322 0.117 ;
        RECT 0.267 0.027 0.285 0.117 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.357 0.099 0.412 0.117 ;
        RECT 0.31 0.063 0.412 0.081 ;
        RECT 0.357 0.063 0.375 0.117 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.171 0.632 0.189 ;
        RECT 0.614 0.063 0.632 0.189 ;
        RECT 0.592 0.063 0.632 0.081 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.445 0.099 0.53 0.117 ;
        RECT 0.512 0.063 0.53 0.117 ;
        RECT 0.445 0.063 0.53 0.081 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.81 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.81 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.702 0.171 0.792 0.189 ;
        RECT 0.774 0.027 0.792 0.189 ;
        RECT 0.701 0.027 0.792 0.045 ;
        RECT 0.702 0.148 0.72 0.189 ;
        RECT 0.701 0.027 0.719 0.068 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.482 0.135 0.567 0.153 ;
      RECT 0.549 0.027 0.567 0.153 ;
      RECT 0.65 0.099 0.695 0.117 ;
      RECT 0.65 0.027 0.668 0.117 ;
      RECT 0.369 0.027 0.668 0.045 ;
      RECT 0.433 0.171 0.549 0.189 ;
      RECT 0.433 0.135 0.451 0.189 ;
      RECT 0.275 0.135 0.451 0.153 ;
      RECT 0.193 0.171 0.392 0.189 ;
      RECT 0.094 0.171 0.135 0.189 ;
    LAYER M2 ;
      RECT 0.099 0.171 0.234 0.189 ;
    LAYER V1 ;
      RECT 0.207 0.171 0.225 0.189 ;
      RECT 0.099 0.171 0.117 0.189 ;
  END
END AO332x2_ASAP7_6t_SL

MACRO AO333x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO333x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.864 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.684 0.135 0.721 0.153 ;
        RECT 0.684 0.063 0.721 0.081 ;
        RECT 0.684 0.063 0.702 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.629 0.063 0.666 0.153 ;
        RECT 0.555 0.099 0.666 0.117 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.027 0.638 0.045 ;
        RECT 0.466 0.063 0.598 0.081 ;
        RECT 0.58 0.027 0.598 0.081 ;
        RECT 0.466 0.099 0.524 0.117 ;
        RECT 0.466 0.063 0.484 0.117 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.205 0.135 0.249 0.153 ;
        RECT 0.231 0.027 0.249 0.153 ;
        RECT 0.202 0.027 0.249 0.045 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.267 0.099 0.322 0.117 ;
        RECT 0.267 0.027 0.322 0.045 ;
        RECT 0.267 0.027 0.285 0.159 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.357 0.099 0.417 0.117 ;
        RECT 0.31 0.063 0.412 0.081 ;
        RECT 0.357 0.063 0.375 0.117 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.159 0.097 0.2 0.115 ;
        RECT 0.159 0.027 0.177 0.158 ;
        RECT 0.094 0.027 0.177 0.045 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.135 0.141 0.153 ;
        RECT 0.123 0.063 0.141 0.153 ;
        RECT 0.093 0.063 0.141 0.081 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.864 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.864 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.796 0.171 0.846 0.189 ;
        RECT 0.828 0.027 0.846 0.189 ;
        RECT 0.796 0.027 0.846 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.634 0.171 0.764 0.189 ;
      RECT 0.746 0.132 0.764 0.189 ;
      RECT 0.757 0.064 0.775 0.152 ;
      RECT 0.746 0.027 0.764 0.084 ;
      RECT 0.688 0.027 0.764 0.045 ;
      RECT 0.585 0.135 0.603 0.176 ;
      RECT 0.313 0.135 0.331 0.176 ;
      RECT 0.313 0.135 0.603 0.153 ;
      RECT 0.505 0.171 0.554 0.189 ;
      RECT 0.364 0.027 0.549 0.045 ;
      RECT 0.363 0.171 0.413 0.189 ;
      RECT 0.193 0.171 0.239 0.189 ;
      RECT 0.094 0.171 0.135 0.189 ;
    LAYER M2 ;
      RECT 0.521 0.171 0.68 0.189 ;
      RECT 0.099 0.171 0.405 0.189 ;
    LAYER V1 ;
      RECT 0.639 0.171 0.657 0.189 ;
      RECT 0.531 0.171 0.549 0.189 ;
      RECT 0.369 0.171 0.387 0.189 ;
      RECT 0.207 0.171 0.225 0.189 ;
      RECT 0.099 0.171 0.117 0.189 ;
  END
END AO333x1_ASAP7_6t_SL

MACRO AO333x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO333x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.918 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.684 0.135 0.721 0.153 ;
        RECT 0.684 0.063 0.721 0.081 ;
        RECT 0.684 0.063 0.702 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.629 0.063 0.666 0.153 ;
        RECT 0.555 0.099 0.666 0.117 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.027 0.638 0.045 ;
        RECT 0.466 0.063 0.598 0.081 ;
        RECT 0.58 0.027 0.598 0.081 ;
        RECT 0.466 0.099 0.522 0.117 ;
        RECT 0.466 0.063 0.484 0.117 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.205 0.135 0.249 0.153 ;
        RECT 0.231 0.027 0.249 0.153 ;
        RECT 0.202 0.027 0.249 0.045 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.267 0.099 0.322 0.117 ;
        RECT 0.267 0.027 0.322 0.045 ;
        RECT 0.267 0.027 0.285 0.159 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.357 0.099 0.412 0.117 ;
        RECT 0.31 0.063 0.412 0.081 ;
        RECT 0.357 0.063 0.375 0.117 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.159 0.097 0.2 0.115 ;
        RECT 0.159 0.027 0.177 0.158 ;
        RECT 0.094 0.027 0.177 0.045 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.135 0.141 0.153 ;
        RECT 0.123 0.063 0.141 0.153 ;
        RECT 0.091 0.063 0.141 0.081 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.063 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.918 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.918 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.796 0.171 0.846 0.189 ;
        RECT 0.828 0.027 0.846 0.189 ;
        RECT 0.796 0.027 0.846 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.634 0.171 0.764 0.189 ;
      RECT 0.746 0.132 0.764 0.189 ;
      RECT 0.757 0.064 0.775 0.152 ;
      RECT 0.746 0.027 0.764 0.084 ;
      RECT 0.688 0.027 0.764 0.045 ;
      RECT 0.585 0.135 0.603 0.176 ;
      RECT 0.313 0.135 0.331 0.176 ;
      RECT 0.313 0.135 0.603 0.153 ;
      RECT 0.505 0.171 0.554 0.189 ;
      RECT 0.364 0.027 0.549 0.045 ;
      RECT 0.363 0.171 0.413 0.189 ;
      RECT 0.193 0.171 0.239 0.189 ;
      RECT 0.094 0.171 0.135 0.189 ;
    LAYER M2 ;
      RECT 0.521 0.171 0.68 0.189 ;
      RECT 0.099 0.171 0.405 0.189 ;
    LAYER V1 ;
      RECT 0.639 0.171 0.657 0.189 ;
      RECT 0.531 0.171 0.549 0.189 ;
      RECT 0.369 0.171 0.387 0.189 ;
      RECT 0.207 0.171 0.225 0.189 ;
      RECT 0.099 0.171 0.117 0.189 ;
  END
END AO333x2_ASAP7_6t_SL

MACRO AO33x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO33x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.187 0.135 0.252 0.153 ;
        RECT 0.234 0.027 0.252 0.153 ;
        RECT 0.202 0.027 0.252 0.064 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.277 0.135 0.317 0.153 ;
        RECT 0.277 0.063 0.315 0.081 ;
        RECT 0.288 0.063 0.306 0.153 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.137 0.099 0.203 0.117 ;
        RECT 0.137 0.027 0.176 0.045 ;
        RECT 0.137 0.027 0.155 0.17 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.34 0.027 0.358 0.11 ;
        RECT 0.28 0.027 0.358 0.045 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.027 0.458 0.045 ;
        RECT 0.376 0.099 0.417 0.117 ;
        RECT 0.376 0.027 0.394 0.117 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.485 0.027 0.524 0.045 ;
        RECT 0.485 0.099 0.522 0.117 ;
        RECT 0.485 0.027 0.503 0.117 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.071 0.135 0.112 0.153 ;
        RECT 0.071 0.055 0.112 0.073 ;
        RECT 0.071 0.027 0.089 0.153 ;
        RECT 0.04 0.027 0.089 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.475 0.171 0.523 0.189 ;
      RECT 0.475 0.135 0.504 0.189 ;
      RECT 0.353 0.135 0.504 0.153 ;
      RECT 0.449 0.063 0.467 0.153 ;
      RECT 0.426 0.063 0.467 0.081 ;
      RECT 0.018 0.171 0.073 0.189 ;
      RECT 0.018 0.092 0.036 0.189 ;
      RECT 0.201 0.171 0.441 0.189 ;
    LAYER M2 ;
      RECT 0.025 0.171 0.514 0.189 ;
    LAYER V1 ;
      RECT 0.477 0.171 0.495 0.189 ;
      RECT 0.045 0.171 0.063 0.189 ;
  END
END AO33x1_ASAP7_6t_SL

MACRO AO33x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO33x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.187 0.135 0.252 0.153 ;
        RECT 0.234 0.027 0.252 0.153 ;
        RECT 0.202 0.027 0.252 0.064 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.277 0.135 0.317 0.153 ;
        RECT 0.277 0.063 0.315 0.081 ;
        RECT 0.288 0.063 0.306 0.153 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.137 0.099 0.203 0.117 ;
        RECT 0.137 0.027 0.176 0.064 ;
        RECT 0.137 0.027 0.155 0.163 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.34 0.027 0.358 0.11 ;
        RECT 0.28 0.027 0.358 0.045 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.027 0.4455 0.045 ;
        RECT 0.376 0.099 0.417 0.117 ;
        RECT 0.376 0.027 0.394 0.117 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.488 0.027 0.531 0.081 ;
        RECT 0.506 0.027 0.524 0.117 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.101 0.104 0.119 0.163 ;
        RECT 0.071 0.055 0.112 0.073 ;
        RECT 0.071 0.104 0.119 0.122 ;
        RECT 0.071 0.027 0.089 0.122 ;
        RECT 0.02 0.027 0.089 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.474 0.171 0.522 0.189 ;
      RECT 0.474 0.135 0.497 0.189 ;
      RECT 0.353 0.135 0.497 0.153 ;
      RECT 0.449 0.063 0.467 0.153 ;
      RECT 0.426 0.063 0.467 0.081 ;
      RECT 0.018 0.17 0.068 0.189 ;
      RECT 0.018 0.092 0.036 0.189 ;
      RECT 0.201 0.171 0.441 0.189 ;
    LAYER M2 ;
      RECT 0.025 0.171 0.513 0.189 ;
    LAYER V1 ;
      RECT 0.477 0.171 0.495 0.189 ;
      RECT 0.045 0.171 0.063 0.189 ;
  END
END AO33x2_ASAP7_6t_SL

MACRO AOI211xp25_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211xp25_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.045 0.144 0.104 ;
        RECT 0.106 0.045 0.144 0.063 ;
      LAYER M2 ;
        RECT 0.063 0.063 0.151 0.081 ;
      LAYER V1 ;
        RECT 0.126 0.063 0.144 0.081 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.07 0.036 0.146 ;
      LAYER M2 ;
        RECT 0.018 0.099 0.098 0.117 ;
      LAYER V1 ;
        RECT 0.018 0.099 0.036 0.117 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.063 0.215 0.081 ;
        RECT 0.178 0.063 0.196 0.122 ;
      LAYER M2 ;
        RECT 0.173 0.099 0.275 0.117 ;
      LAYER V1 ;
        RECT 0.178 0.099 0.196 0.117 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.217 0.135 0.254 0.153 ;
        RECT 0.236 0.094 0.254 0.153 ;
      LAYER M2 ;
        RECT 0.159 0.135 0.243 0.153 ;
      LAYER V1 ;
        RECT 0.22 0.135 0.238 0.153 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.247 0.171 0.306 0.189 ;
        RECT 0.288 0.027 0.306 0.189 ;
        RECT 0.18 0.027 0.306 0.045 ;
        RECT 0.063 0.135 0.117 0.153 ;
        RECT 0.063 0.027 0.081 0.153 ;
        RECT 0.04 0.027 0.081 0.045 ;
      LAYER M2 ;
        RECT 0.04 0.027 0.279 0.045 ;
      LAYER V1 ;
        RECT 0.045 0.027 0.063 0.045 ;
        RECT 0.261 0.027 0.279 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.171 0.176 0.189 ;
  END
END AOI211xp25_ASAP7_6t_SL

MACRO AOI211xp5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211xp5_ASAP7_6t_SL 0 0 ;
  SIZE 0.648 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.118 0.117 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.648 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.177 0.099 0.245 0.117 ;
      LAYER M1 ;
        RECT 0.159 0.099 0.238 0.117 ;
        RECT 0.159 0.135 0.234 0.153 ;
        RECT 0.159 0.027 0.234 0.045 ;
        RECT 0.159 0.027 0.177 0.153 ;
      LAYER V1 ;
        RECT 0.202 0.099 0.22 0.117 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.289 0.063 0.357 0.081 ;
      LAYER M1 ;
        RECT 0.314 0.099 0.369 0.117 ;
        RECT 0.314 0.027 0.369 0.045 ;
        RECT 0.314 0.027 0.332 0.117 ;
      LAYER V1 ;
        RECT 0.314 0.063 0.332 0.081 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.495 0.099 0.563 0.117 ;
      LAYER M1 ;
        RECT 0.512 0.099 0.567 0.117 ;
        RECT 0.549 0.063 0.567 0.117 ;
        RECT 0.512 0.063 0.567 0.081 ;
      LAYER V1 ;
        RECT 0.52 0.099 0.538 0.117 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.094 0.027 0.608 0.045 ;
      LAYER M1 ;
        RECT 0.519 0.135 0.637 0.153 ;
        RECT 0.619 0.027 0.637 0.153 ;
        RECT 0.583 0.027 0.637 0.045 ;
        RECT 0.453 0.027 0.5 0.045 ;
        RECT 0.094 0.027 0.131 0.045 ;
      LAYER V1 ;
        RECT 0.099 0.027 0.117 0.045 ;
        RECT 0.477 0.027 0.495 0.045 ;
        RECT 0.585 0.027 0.603 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.171 0.306 0.189 ;
      RECT 0.288 0.135 0.306 0.189 ;
      RECT 0.288 0.135 0.449 0.153 ;
      RECT 0.361 0.171 0.608 0.189 ;
  END
END AOI211xp5_ASAP7_6t_SL

MACRO AOI21x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.158 0.099 0.333 0.117 ;
        RECT 0.139 0.135 0.176 0.153 ;
        RECT 0.158 0.063 0.176 0.153 ;
        RECT 0.139 0.063 0.176 0.081 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.098 0.077 0.116 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.364 0.099 0.461 0.117 ;
        RECT 0.443 0.063 0.461 0.117 ;
        RECT 0.395 0.063 0.461 0.081 ;
        RECT 0.305 0.135 0.382 0.153 ;
        RECT 0.364 0.099 0.382 0.153 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.418 0.135 0.514 0.153 ;
        RECT 0.496 0.027 0.514 0.153 ;
        RECT 0.256 0.027 0.514 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.207 0.063 0.338 0.081 ;
      RECT 0.207 0.027 0.225 0.081 ;
      RECT 0.094 0.027 0.225 0.045 ;
      RECT 0.094 0.171 0.5 0.189 ;
  END
END AOI21x1_ASAP7_6t_SL

MACRO AOI21xp25_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21xp25_ASAP7_6t_SL 0 0 ;
  SIZE 0.27 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.086 0.098 0.146 0.116 ;
        RECT 0.086 0.027 0.123 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.028 0.116 0.068 0.153 ;
        RECT 0.028 0.027 0.068 0.072 ;
        RECT 0.028 0.027 0.046 0.153 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.135 0.217 0.153 ;
        RECT 0.18 0.063 0.217 0.081 ;
        RECT 0.18 0.063 0.198 0.153 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.27 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.27 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.171 0.261 0.189 ;
        RECT 0.243 0.027 0.261 0.189 ;
        RECT 0.148 0.027 0.261 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.171 0.171 0.189 ;
  END
END AOI21xp25_ASAP7_6t_SL

MACRO AOI21xp5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21xp5_ASAP7_6t_SL 0 0 ;
  SIZE 0.27 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.086 0.098 0.146 0.116 ;
        RECT 0.086 0.027 0.123 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.028 0.116 0.068 0.153 ;
        RECT 0.028 0.027 0.068 0.068 ;
        RECT 0.028 0.027 0.046 0.153 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.135 0.217 0.153 ;
        RECT 0.18 0.063 0.217 0.081 ;
        RECT 0.18 0.063 0.198 0.153 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.27 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.27 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.171 0.261 0.189 ;
        RECT 0.243 0.027 0.261 0.189 ;
        RECT 0.148 0.027 0.261 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.171 0.171 0.189 ;
  END
END AOI21xp5_ASAP7_6t_SL

MACRO AOI221xp25_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221xp25_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.238 0.135 0.293 0.153 ;
        RECT 0.275 0.027 0.293 0.153 ;
        RECT 0.234 0.099 0.293 0.117 ;
        RECT 0.256 0.027 0.293 0.045 ;
      LAYER M2 ;
        RECT 0.217 0.135 0.309 0.153 ;
      LAYER V1 ;
        RECT 0.252 0.135 0.27 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.311 0.116 0.36 0.153 ;
        RECT 0.342 0.028 0.36 0.153 ;
        RECT 0.311 0.028 0.36 0.065 ;
      LAYER M2 ;
        RECT 0.296 0.099 0.36 0.117 ;
      LAYER V1 ;
        RECT 0.342 0.099 0.36 0.117 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.058 0.036 0.151 ;
      LAYER M2 ;
        RECT 0.018 0.099 0.082 0.117 ;
      LAYER V1 ;
        RECT 0.018 0.099 0.036 0.117 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.063 0.144 0.11 ;
        RECT 0.106 0.063 0.144 0.081 ;
      LAYER M2 ;
        RECT 0.097 0.063 0.161 0.081 ;
      LAYER V1 ;
        RECT 0.113 0.063 0.131 0.081 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.063 0.217 0.081 ;
        RECT 0.16 0.135 0.198 0.153 ;
        RECT 0.18 0.063 0.198 0.153 ;
      LAYER M2 ;
        RECT 0.157 0.099 0.221 0.117 ;
      LAYER V1 ;
        RECT 0.18 0.099 0.198 0.117 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.063 0.027 0.225 0.045 ;
        RECT 0.063 0.135 0.122 0.153 ;
        RECT 0.063 0.027 0.081 0.153 ;
      LAYER M2 ;
        RECT 0.0495 0.135 0.12 0.153 ;
      LAYER V1 ;
        RECT 0.078 0.135 0.096 0.153 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.207 0.171 0.338 0.189 ;
      RECT 0.04 0.171 0.176 0.189 ;
  END
END AOI221xp25_ASAP7_6t_SL

MACRO AOI221xp5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221xp5_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.254 0.063 0.292 0.081 ;
        RECT 0.254 0.135 0.291 0.153 ;
        RECT 0.254 0.063 0.272 0.153 ;
        RECT 0.231 0.096 0.272 0.114 ;
      LAYER M2 ;
        RECT 0.178 0.063 0.282 0.081 ;
      LAYER V1 ;
        RECT 0.259 0.063 0.277 0.081 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.323 0.116 0.362 0.153 ;
        RECT 0.344 0.027 0.362 0.153 ;
        RECT 0.309 0.027 0.362 0.045 ;
      LAYER M2 ;
        RECT 0.258 0.099 0.362 0.117 ;
      LAYER V1 ;
        RECT 0.344 0.099 0.362 0.117 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.053 0.047 0.09 ;
        RECT 0.018 0.053 0.036 0.122 ;
      LAYER M2 ;
        RECT 0.024 0.063 0.128 0.081 ;
      LAYER V1 ;
        RECT 0.029 0.063 0.047 0.081 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.129 0.063 0.147 0.119 ;
        RECT 0.108 0.063 0.147 0.081 ;
      LAYER M2 ;
        RECT 0.045 0.099 0.147 0.117 ;
      LAYER V1 ;
        RECT 0.129 0.099 0.147 0.117 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.159 0.135 0.223 0.153 ;
        RECT 0.172 0.063 0.214 0.081 ;
        RECT 0.18 0.063 0.198 0.153 ;
      LAYER M2 ;
        RECT 0.169 0.135 0.273 0.153 ;
      LAYER V1 ;
        RECT 0.174 0.135 0.192 0.153 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.065 0.027 0.225 0.045 ;
        RECT 0.065 0.135 0.112 0.153 ;
        RECT 0.065 0.027 0.083 0.153 ;
      LAYER M2 ;
        RECT 0.047 0.027 0.204 0.045 ;
      LAYER V1 ;
        RECT 0.099 0.027 0.117 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.202 0.171 0.338 0.189 ;
      RECT 0.04 0.171 0.171 0.189 ;
  END
END AOI221xp5_ASAP7_6t_SL

MACRO AOI222xp25_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222xp25_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.058 0.036 0.146 ;
      LAYER M2 ;
        RECT 0.018 0.099 0.088 0.117 ;
      LAYER V1 ;
        RECT 0.018 0.099 0.036 0.117 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.063 0.144 0.117 ;
        RECT 0.106 0.063 0.144 0.081 ;
      LAYER M2 ;
        RECT 0.103 0.063 0.187 0.081 ;
      LAYER V1 ;
        RECT 0.112 0.063 0.13 0.081 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.099 0.355 0.117 ;
        RECT 0.337 0.063 0.355 0.117 ;
        RECT 0.3 0.063 0.355 0.081 ;
      LAYER M2 ;
        RECT 0.287 0.063 0.371 0.081 ;
      LAYER V1 ;
        RECT 0.313 0.063 0.331 0.081 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.182 0.099 0.237 0.117 ;
        RECT 0.182 0.063 0.237 0.081 ;
        RECT 0.182 0.063 0.2 0.117 ;
      LAYER M2 ;
        RECT 0.164 0.099 0.238 0.117 ;
      LAYER V1 ;
        RECT 0.2 0.099 0.218 0.117 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.416 0.116 0.453 0.153 ;
        RECT 0.416 0.027 0.453 0.064 ;
        RECT 0.416 0.027 0.434 0.153 ;
        RECT 0.393 0.097 0.434 0.115 ;
      LAYER M2 ;
        RECT 0.361 0.099 0.46 0.117 ;
      LAYER V1 ;
        RECT 0.416 0.099 0.434 0.117 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.471 0.15 0.524 0.189 ;
        RECT 0.506 0.027 0.524 0.189 ;
        RECT 0.472 0.027 0.524 0.064 ;
      LAYER M2 ;
        RECT 0.447 0.171 0.524 0.189 ;
      LAYER V1 ;
        RECT 0.477 0.171 0.495 0.189 ;
    END
  END C2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.063 0.027 0.338 0.045 ;
        RECT 0.063 0.135 0.117 0.153 ;
        RECT 0.063 0.027 0.081 0.153 ;
      LAYER M2 ;
        RECT 0.055 0.135 0.132 0.153 ;
      LAYER V1 ;
        RECT 0.082 0.135 0.1 0.153 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.342 0.171 0.446 0.189 ;
      RECT 0.342 0.135 0.36 0.189 ;
      RECT 0.199 0.135 0.36 0.153 ;
      RECT 0.04 0.171 0.284 0.189 ;
  END
END AOI222xp25_ASAP7_6t_SL

MACRO AOI22xp25_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22xp25_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.031 0.116 0.068 0.153 ;
        RECT 0.031 0.027 0.068 0.064 ;
        RECT 0.031 0.027 0.049 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.105 0.098 0.141 0.116 ;
        RECT 0.086 0.116 0.123 0.153 ;
        RECT 0.105 0.027 0.123 0.153 ;
        RECT 0.086 0.027 0.123 0.064 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.116 0.294 0.153 ;
        RECT 0.276 0.027 0.294 0.153 ;
        RECT 0.256 0.027 0.294 0.045 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.135 0.191 0.153 ;
        RECT 0.173 0.027 0.191 0.153 ;
        RECT 0.141 0.027 0.191 0.064 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.211 0.055 0.229 0.158 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.248 0.171 0.285 0.189 ;
      RECT 0.04 0.171 0.176 0.189 ;
    LAYER M2 ;
      RECT 0.148 0.171 0.284 0.189 ;
    LAYER V1 ;
      RECT 0.261 0.171 0.279 0.189 ;
      RECT 0.153 0.171 0.171 0.189 ;
  END
END AOI22xp25_ASAP7_6t_SL

MACRO AOI22xp5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22xp5_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.031 0.116 0.068 0.153 ;
        RECT 0.031 0.027 0.068 0.064 ;
        RECT 0.031 0.027 0.049 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.105 0.098 0.141 0.116 ;
        RECT 0.086 0.116 0.123 0.153 ;
        RECT 0.105 0.027 0.123 0.153 ;
        RECT 0.086 0.027 0.123 0.064 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.116 0.294 0.153 ;
        RECT 0.276 0.027 0.294 0.153 ;
        RECT 0.256 0.027 0.294 0.045 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.135 0.191 0.153 ;
        RECT 0.173 0.027 0.191 0.153 ;
        RECT 0.141 0.027 0.191 0.064 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.211 0.055 0.229 0.158 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.248 0.171 0.285 0.189 ;
      RECT 0.04 0.171 0.176 0.189 ;
    LAYER M2 ;
      RECT 0.148 0.171 0.284 0.189 ;
    LAYER V1 ;
      RECT 0.261 0.171 0.279 0.189 ;
      RECT 0.153 0.171 0.171 0.189 ;
  END
END AOI22xp5_ASAP7_6t_SL

MACRO AOI311xp33_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI311xp33_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.17 0.063 0.207 0.081 ;
        RECT 0.18 0.063 0.198 0.122 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.135 0.144 0.153 ;
        RECT 0.126 0.027 0.144 0.153 ;
        RECT 0.094 0.027 0.144 0.045 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.09 0.117 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.215 0.135 0.252 0.153 ;
        RECT 0.234 0.094 0.252 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.277 0.135 0.317 0.153 ;
        RECT 0.28 0.063 0.317 0.081 ;
        RECT 0.288 0.063 0.306 0.153 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.302 0.171 0.36 0.189 ;
        RECT 0.342 0.027 0.36 0.189 ;
        RECT 0.198 0.027 0.36 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.171 0.234 0.189 ;
  END
END AOI311xp33_ASAP7_6t_SL

MACRO AOI31xp33_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31xp33_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.159 0.116 0.204 0.153 ;
        RECT 0.177 0.064 0.195 0.153 ;
        RECT 0.166 0.064 0.195 0.082 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.116 0.141 0.153 ;
        RECT 0.123 0.027 0.141 0.153 ;
        RECT 0.091 0.027 0.141 0.064 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.152 0.069 0.189 ;
        RECT 0.017 0.027 0.068 0.064 ;
        RECT 0.017 0.027 0.035 0.189 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.227 0.063 0.265 0.083 ;
        RECT 0.225 0.116 0.262 0.153 ;
        RECT 0.234 0.063 0.252 0.153 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.29 0.027 0.308 0.182 ;
        RECT 0.202 0.027 0.308 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.171 0.23 0.189 ;
  END
END AOI31xp33_ASAP7_6t_SL

MACRO AOI31xp67_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31xp67_ASAP7_6t_SL 0 0 ;
  SIZE 0.702 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.513 0.099 0.689 0.117 ;
        RECT 0.671 0.063 0.689 0.117 ;
        RECT 0.634 0.063 0.689 0.081 ;
        RECT 0.58 0.171 0.617 0.189 ;
        RECT 0.58 0.099 0.598 0.189 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.273 0.099 0.466 0.117 ;
        RECT 0.273 0.135 0.328 0.153 ;
        RECT 0.273 0.027 0.328 0.045 ;
        RECT 0.273 0.027 0.291 0.153 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.095 0.117 ;
        RECT 0.018 0.135 0.073 0.153 ;
        RECT 0.018 0.027 0.063 0.045 ;
        RECT 0.018 0.027 0.036 0.153 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.154 0.098 0.209 0.116 ;
        RECT 0.121 0.135 0.172 0.153 ;
        RECT 0.154 0.063 0.172 0.153 ;
        RECT 0.117 0.063 0.172 0.081 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.702 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.702 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.207 0.135 0.663 0.153 ;
      LAYER M1 ;
        RECT 0.629 0.135 0.674 0.153 ;
        RECT 0.2 0.135 0.255 0.153 ;
        RECT 0.237 0.027 0.255 0.153 ;
        RECT 0.202 0.027 0.255 0.045 ;
      LAYER V1 ;
        RECT 0.232 0.135 0.25 0.153 ;
        RECT 0.64 0.135 0.658 0.153 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.526 0.027 0.663 0.045 ;
      RECT 0.364 0.063 0.603 0.081 ;
      RECT 0.04 0.171 0.554 0.189 ;
      RECT 0.408 0.027 0.447 0.045 ;
      RECT 0.094 0.027 0.131 0.045 ;
    LAYER M2 ;
      RECT 0.094 0.027 0.447 0.045 ;
    LAYER V1 ;
      RECT 0.423 0.027 0.441 0.045 ;
      RECT 0.099 0.027 0.117 0.045 ;
  END
END AOI31xp67_ASAP7_6t_SL

MACRO AOI321xp17_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI321xp17_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.07 0.198 0.122 ;
      LAYER M2 ;
        RECT 0.158 0.099 0.222 0.117 ;
      LAYER V1 ;
        RECT 0.18 0.099 0.198 0.117 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.135 0.144 0.153 ;
        RECT 0.126 0.027 0.144 0.153 ;
        RECT 0.094 0.027 0.144 0.045 ;
      LAYER M2 ;
        RECT 0.097 0.135 0.163 0.153 ;
      LAYER V1 ;
        RECT 0.124 0.135 0.142 0.153 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
      LAYER M2 ;
        RECT 0.018 0.099 0.106 0.117 ;
      LAYER V1 ;
        RECT 0.018 0.099 0.036 0.117 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.277 0.027 0.317 0.045 ;
        RECT 0.285 0.027 0.303 0.119 ;
      LAYER M2 ;
        RECT 0.257 0.099 0.321 0.117 ;
      LAYER V1 ;
        RECT 0.285 0.099 0.303 0.117 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.36 0.063 0.378 0.11 ;
        RECT 0.341 0.063 0.378 0.081 ;
      LAYER M2 ;
        RECT 0.339 0.063 0.403 0.081 ;
      LAYER V1 ;
        RECT 0.351 0.063 0.369 0.081 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.135 0.271 0.153 ;
        RECT 0.234 0.07 0.252 0.153 ;
      LAYER M2 ;
        RECT 0.212 0.135 0.278 0.153 ;
      LAYER V1 ;
        RECT 0.236 0.135 0.254 0.153 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.315 0.135 0.414 0.153 ;
        RECT 0.396 0.027 0.414 0.153 ;
        RECT 0.356 0.027 0.414 0.045 ;
        RECT 0.198 0.027 0.238 0.045 ;
      LAYER M2 ;
        RECT 0.207 0.027 0.392 0.045 ;
      LAYER V1 ;
        RECT 0.207 0.027 0.225 0.045 ;
        RECT 0.369 0.027 0.387 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.256 0.171 0.396 0.189 ;
      RECT 0.094 0.171 0.225 0.189 ;
  END
END AOI321xp17_ASAP7_6t_SL

MACRO AOI322xp17_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI322xp17_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.135 0.071 0.153 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.153 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.141 0.099 0.22 0.117 ;
      LAYER M1 ;
        RECT 0.159 0.099 0.196 0.117 ;
        RECT 0.159 0.061 0.177 0.117 ;
      LAYER V1 ;
        RECT 0.17 0.099 0.188 0.117 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.202 0.063 0.27 0.081 ;
      LAYER M1 ;
        RECT 0.234 0.063 0.252 0.11 ;
        RECT 0.205 0.063 0.252 0.081 ;
      LAYER V1 ;
        RECT 0.207 0.063 0.225 0.081 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.271 0.135 0.362 0.153 ;
      LAYER M1 ;
        RECT 0.292 0.135 0.333 0.153 ;
        RECT 0.28 0.027 0.317 0.045 ;
        RECT 0.292 0.088 0.31 0.153 ;
        RECT 0.288 0.027 0.306 0.106 ;
      LAYER V1 ;
        RECT 0.302 0.135 0.32 0.153 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.076 0.063 0.153 0.081 ;
      LAYER M1 ;
        RECT 0.084 0.099 0.141 0.117 ;
        RECT 0.123 0.027 0.141 0.117 ;
        RECT 0.094 0.027 0.141 0.045 ;
      LAYER V1 ;
        RECT 0.123 0.063 0.141 0.081 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.378 0.063 0.448 0.081 ;
      LAYER M1 ;
        RECT 0.412 0.063 0.43 0.11 ;
        RECT 0.388 0.063 0.43 0.081 ;
      LAYER V1 ;
        RECT 0.39 0.063 0.408 0.081 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.326 0.099 0.4 0.117 ;
      LAYER M1 ;
        RECT 0.342 0.099 0.379 0.117 ;
        RECT 0.342 0.027 0.379 0.045 ;
        RECT 0.342 0.027 0.36 0.117 ;
      LAYER V1 ;
        RECT 0.351 0.099 0.369 0.117 ;
    END
  END C2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.202 0.027 0.446 0.045 ;
      LAYER M1 ;
        RECT 0.364 0.135 0.468 0.153 ;
        RECT 0.45 0.027 0.468 0.153 ;
        RECT 0.413 0.027 0.468 0.045 ;
        RECT 0.194 0.027 0.249 0.045 ;
      LAYER V1 ;
        RECT 0.207 0.027 0.225 0.045 ;
        RECT 0.423 0.027 0.441 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.171 0.176 0.189 ;
      RECT 0.102 0.135 0.12 0.189 ;
      RECT 0.102 0.135 0.267 0.153 ;
      RECT 0.207 0.171 0.45 0.189 ;
  END
END AOI322xp17_ASAP7_6t_SL

MACRO AOI32xp33_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32xp33_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.016 0.027 0.068 0.045 ;
        RECT 0.016 0.027 0.034 0.127 ;
      LAYER M2 ;
        RECT 0.038 0.027 0.168 0.045 ;
      LAYER V1 ;
        RECT 0.045 0.027 0.063 0.045 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.078 0.099 0.149 0.117 ;
      LAYER M2 ;
        RECT 0.061 0.099 0.163 0.117 ;
      LAYER V1 ;
        RECT 0.1 0.099 0.118 0.117 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.135 0.221 0.153 ;
        RECT 0.18 0.088 0.198 0.153 ;
      LAYER M2 ;
        RECT 0.147 0.135 0.249 0.153 ;
      LAYER V1 ;
        RECT 0.193 0.135 0.211 0.153 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.232 0.063 0.27 0.081 ;
        RECT 0.232 0.063 0.25 0.118 ;
      LAYER M2 ;
        RECT 0.215 0.063 0.307 0.081 ;
      LAYER V1 ;
        RECT 0.249 0.063 0.267 0.081 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.279 0.099 0.327 0.117 ;
        RECT 0.309 0.07 0.327 0.117 ;
      LAYER M2 ;
        RECT 0.243 0.099 0.345 0.117 ;
      LAYER V1 ;
        RECT 0.284 0.099 0.302 0.117 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.135 0.363 0.153 ;
        RECT 0.345 0.027 0.363 0.153 ;
        RECT 0.148 0.027 0.363 0.045 ;
        RECT 0.261 0.135 0.279 0.176 ;
      LAYER M2 ;
        RECT 0.209 0.027 0.338 0.045 ;
      LAYER V1 ;
        RECT 0.315 0.027 0.333 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.31 0.171 0.347 0.189 ;
      RECT 0.094 0.171 0.23 0.189 ;
    LAYER M2 ;
      RECT 0.148 0.171 0.338 0.189 ;
    LAYER V1 ;
      RECT 0.315 0.171 0.333 0.189 ;
      RECT 0.153 0.171 0.171 0.189 ;
  END
END AOI32xp33_ASAP7_6t_SL

MACRO AOI331xp17_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI331xp17_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.135 0.224 0.153 ;
        RECT 0.18 0.07 0.198 0.153 ;
      LAYER M2 ;
        RECT 0.182 0.135 0.272 0.153 ;
      LAYER V1 ;
        RECT 0.2 0.135 0.218 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.135 0.155 0.153 ;
        RECT 0.094 0.027 0.155 0.045 ;
        RECT 0.126 0.027 0.144 0.153 ;
      LAYER M2 ;
        RECT 0.0885 0.063 0.1775 0.081 ;
      LAYER V1 ;
        RECT 0.126 0.063 0.144 0.081 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.171 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
      LAYER M2 ;
        RECT 0.038 0.171 0.136 0.189 ;
      LAYER V1 ;
        RECT 0.045 0.171 0.063 0.189 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.099 0.271 0.117 ;
        RECT 0.234 0.07 0.252 0.117 ;
      LAYER M2 ;
        RECT 0.172 0.099 0.298 0.117 ;
      LAYER V1 ;
        RECT 0.237 0.099 0.255 0.117 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.278 0.027 0.315 0.045 ;
        RECT 0.288 0.027 0.306 0.088 ;
      LAYER M2 ;
        RECT 0.212 0.063 0.311 0.081 ;
      LAYER V1 ;
        RECT 0.288 0.063 0.306 0.081 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.027 0.379 0.045 ;
        RECT 0.342 0.027 0.36 0.108 ;
      LAYER M2 ;
        RECT 0.342 0.063 0.42 0.081 ;
      LAYER V1 ;
        RECT 0.342 0.063 0.36 0.081 ;
    END
  END B3
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.412 0.07 0.43 0.14 ;
      LAYER M2 ;
        RECT 0.364 0.099 0.453 0.117 ;
      LAYER V1 ;
        RECT 0.412 0.099 0.43 0.117 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.418 0.171 0.468 0.189 ;
        RECT 0.45 0.027 0.468 0.189 ;
        RECT 0.41 0.027 0.468 0.045 ;
        RECT 0.195 0.027 0.237 0.045 ;
      LAYER M2 ;
        RECT 0.201 0.027 0.451 0.045 ;
      LAYER V1 ;
        RECT 0.207 0.027 0.225 0.045 ;
        RECT 0.423 0.027 0.441 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.369 0.135 0.387 0.181 ;
      RECT 0.256 0.135 0.387 0.153 ;
      RECT 0.099 0.171 0.338 0.189 ;
  END
END AOI331xp17_ASAP7_6t_SL

MACRO AOI332xp17_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI332xp17_ASAP7_6t_SL 0 0 ;
  SIZE 0.594 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.159 0.097 0.201 0.115 ;
        RECT 0.159 0.027 0.177 0.158 ;
        RECT 0.094 0.027 0.177 0.045 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.135 0.141 0.153 ;
        RECT 0.123 0.063 0.141 0.153 ;
        RECT 0.08 0.063 0.141 0.081 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.063 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.135 0.249 0.153 ;
        RECT 0.231 0.027 0.249 0.153 ;
        RECT 0.202 0.027 0.249 0.045 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.267 0.027 0.333 0.045 ;
        RECT 0.267 0.099 0.322 0.117 ;
        RECT 0.267 0.027 0.285 0.117 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.357 0.099 0.416 0.117 ;
        RECT 0.31 0.063 0.412 0.081 ;
        RECT 0.357 0.063 0.375 0.117 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.557 0.051 0.575 0.14 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.448 0.099 0.503 0.117 ;
        RECT 0.485 0.063 0.503 0.117 ;
        RECT 0.445 0.063 0.503 0.081 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.594 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.482 0.135 0.539 0.153 ;
        RECT 0.521 0.027 0.539 0.153 ;
        RECT 0.364 0.027 0.539 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.433 0.171 0.568 0.189 ;
      RECT 0.433 0.135 0.451 0.189 ;
      RECT 0.275 0.135 0.451 0.153 ;
      RECT 0.201 0.171 0.392 0.189 ;
      RECT 0.094 0.171 0.135 0.189 ;
    LAYER M2 ;
      RECT 0.099 0.171 0.234 0.189 ;
    LAYER V1 ;
      RECT 0.207 0.171 0.225 0.189 ;
      RECT 0.099 0.171 0.117 0.189 ;
  END
END AOI332xp17_ASAP7_6t_SL

MACRO AOI333xp17_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI333xp17_ASAP7_6t_SL 0 0 ;
  SIZE 0.702 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.027 0.662 0.045 ;
        RECT 0.638 0.027 0.656 0.129 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.559 0.099 0.617 0.117 ;
        RECT 0.599 0.063 0.617 0.117 ;
        RECT 0.559 0.063 0.617 0.081 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.464 0.099 0.522 0.117 ;
        RECT 0.464 0.063 0.521 0.081 ;
        RECT 0.464 0.063 0.482 0.117 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.027 0.284 0.045 ;
        RECT 0.237 0.027 0.255 0.116 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.291 0.099 0.36 0.117 ;
        RECT 0.342 0.063 0.36 0.117 ;
        RECT 0.295 0.063 0.36 0.081 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.389 0.099 0.446 0.117 ;
        RECT 0.428 0.063 0.446 0.117 ;
        RECT 0.391 0.063 0.446 0.081 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.135 0.23 0.153 ;
        RECT 0.178 0.067 0.196 0.153 ;
        RECT 0.159 0.067 0.196 0.088 ;
        RECT 0.159 0.027 0.177 0.088 ;
        RECT 0.105 0.027 0.177 0.045 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.086 0.135 0.141 0.153 ;
        RECT 0.123 0.063 0.141 0.153 ;
        RECT 0.08 0.063 0.141 0.081 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.07 0.045 ;
        RECT 0.018 0.027 0.036 0.163 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.702 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.702 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.521 0.171 0.68 0.189 ;
      LAYER M1 ;
        RECT 0.633 0.171 0.692 0.189 ;
        RECT 0.674 0.064 0.692 0.189 ;
        RECT 0.505 0.171 0.554 0.189 ;
      LAYER V1 ;
        RECT 0.531 0.171 0.549 0.189 ;
        RECT 0.639 0.171 0.657 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.585 0.135 0.603 0.176 ;
      RECT 0.265 0.135 0.283 0.176 ;
      RECT 0.265 0.135 0.603 0.153 ;
      RECT 0.315 0.027 0.549 0.045 ;
      RECT 0.315 0.171 0.393 0.189 ;
      RECT 0.187 0.171 0.23 0.189 ;
      RECT 0.086 0.171 0.135 0.189 ;
    LAYER M2 ;
      RECT 0.094 0.171 0.393 0.189 ;
    LAYER V1 ;
      RECT 0.369 0.171 0.387 0.189 ;
      RECT 0.207 0.171 0.225 0.189 ;
      RECT 0.099 0.171 0.117 0.189 ;
  END
END AOI333xp17_ASAP7_6t_SL

MACRO AOI33xp33_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33xp33_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.171 0.055 0.189 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.086 0.099 0.142 0.117 ;
        RECT 0.086 0.027 0.123 0.045 ;
        RECT 0.065 0.135 0.104 0.153 ;
        RECT 0.086 0.027 0.104 0.153 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.161 0.135 0.198 0.153 ;
        RECT 0.18 0.063 0.198 0.153 ;
        RECT 0.134 0.063 0.198 0.081 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.252 0.027 0.312 0.045 ;
        RECT 0.252 0.099 0.289 0.117 ;
        RECT 0.252 0.027 0.27 0.117 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.321 0.099 0.381 0.117 ;
        RECT 0.363 0.027 0.381 0.117 ;
        RECT 0.344 0.027 0.381 0.045 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.459 0.027 0.477 0.165 ;
        RECT 0.412 0.099 0.477 0.117 ;
        RECT 0.44 0.027 0.477 0.045 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.423 0.135 0.441 0.176 ;
        RECT 0.216 0.135 0.441 0.153 ;
        RECT 0.216 0.027 0.234 0.153 ;
        RECT 0.176 0.027 0.234 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.086 0.171 0.392 0.189 ;
  END
END AOI33xp33_ASAP7_6t_SL

MACRO BUFx10_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx10_ASAP7_6t_SL 0 0 ;
  SIZE 0.756 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.095 0.117 ;
        RECT 0.018 0.171 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.756 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.756 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.171 0.738 0.189 ;
        RECT 0.72 0.027 0.738 0.189 ;
        RECT 0.202 0.027 0.738 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.099 0.171 0.144 0.189 ;
      RECT 0.126 0.027 0.144 0.189 ;
      RECT 0.126 0.099 0.689 0.117 ;
      RECT 0.099 0.027 0.144 0.045 ;
  END
END BUFx10_ASAP7_6t_SL

MACRO BUFx12_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx12_ASAP7_6t_SL 0 0 ;
  SIZE 0.864 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.864 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.864 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.171 0.846 0.189 ;
        RECT 0.828 0.027 0.846 0.189 ;
        RECT 0.202 0.027 0.846 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.171 0.144 0.189 ;
      RECT 0.126 0.027 0.144 0.189 ;
      RECT 0.126 0.099 0.797 0.117 ;
      RECT 0.094 0.027 0.144 0.045 ;
  END
END BUFx12_ASAP7_6t_SL

MACRO BUFx12q_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx12q_ASAP7_6t_SL 0 0 ;
  SIZE 0.972 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.02 0.099 0.095 0.117 ;
        RECT 0.02 0.152 0.068 0.189 ;
        RECT 0.02 0.027 0.068 0.064 ;
        RECT 0.02 0.027 0.038 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.972 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.972 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.31 0.171 0.954 0.189 ;
        RECT 0.936 0.027 0.954 0.189 ;
        RECT 0.31 0.027 0.954 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.171 0.279 0.189 ;
      RECT 0.261 0.027 0.279 0.189 ;
      RECT 0.261 0.099 0.311 0.117 ;
      RECT 0.094 0.027 0.279 0.045 ;
  END
END BUFx12q_ASAP7_6t_SL

MACRO BUFx16q_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx16q_ASAP7_6t_SL 0 0 ;
  SIZE 1.188 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.099 0.095 0.117 ;
        RECT 0.017 0.152 0.068 0.189 ;
        RECT 0.017 0.027 0.068 0.064 ;
        RECT 0.017 0.027 0.035 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.188 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.188 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.31 0.171 1.17 0.189 ;
        RECT 1.152 0.027 1.17 0.189 ;
        RECT 0.31 0.027 1.17 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.171 0.252 0.189 ;
      RECT 0.234 0.027 0.252 0.189 ;
      RECT 0.234 0.099 1.121 0.117 ;
      RECT 0.094 0.027 0.252 0.045 ;
  END
END BUFx16q_ASAP7_6t_SL

MACRO BUFx24_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx24_ASAP7_6t_SL 0 0 ;
  SIZE 1.62 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.186 0.117 ;
        RECT 0.018 0.171 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.62 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.62 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.31 0.171 1.602 0.189 ;
        RECT 1.584 0.027 1.602 0.189 ;
        RECT 0.31 0.027 1.602 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.099 0.171 0.252 0.189 ;
      RECT 0.234 0.027 0.252 0.189 ;
      RECT 0.234 0.099 1.553 0.117 ;
      RECT 0.099 0.027 0.252 0.045 ;
  END
END BUFx24_ASAP7_6t_SL

MACRO BUFx2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx2_ASAP7_6t_SL 0 0 ;
  SIZE 0.27 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.078 0.117 ;
        RECT 0.018 0.135 0.073 0.153 ;
        RECT 0.018 0.063 0.073 0.081 ;
        RECT 0.018 0.063 0.036 0.153 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.27 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.27 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.171 0.252 0.189 ;
        RECT 0.234 0.027 0.252 0.189 ;
        RECT 0.148 0.027 0.252 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.171 0.122 0.189 ;
      RECT 0.104 0.027 0.122 0.189 ;
      RECT 0.104 0.099 0.203 0.117 ;
      RECT 0.04 0.027 0.122 0.045 ;
  END
END BUFx2_ASAP7_6t_SL

MACRO BUFx3_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx3_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.01 0.099 0.078 0.117 ;
        RECT 0.01 0.135 0.074 0.153 ;
        RECT 0.01 0.063 0.074 0.081 ;
        RECT 0.01 0.063 0.028 0.153 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.171 0.306 0.189 ;
        RECT 0.288 0.027 0.306 0.189 ;
        RECT 0.148 0.027 0.306 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.171 0.122 0.189 ;
      RECT 0.104 0.027 0.122 0.189 ;
      RECT 0.104 0.099 0.257 0.117 ;
      RECT 0.04 0.027 0.122 0.045 ;
  END
END BUFx3_ASAP7_6t_SL

MACRO BUFx4_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx4_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.01 0.099 0.078 0.117 ;
        RECT 0.01 0.135 0.068 0.153 ;
        RECT 0.01 0.063 0.068 0.081 ;
        RECT 0.01 0.063 0.028 0.153 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.171 0.357 0.189 ;
        RECT 0.339 0.027 0.357 0.189 ;
        RECT 0.148 0.027 0.357 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.171 0.122 0.189 ;
      RECT 0.104 0.027 0.122 0.189 ;
      RECT 0.104 0.099 0.311 0.117 ;
      RECT 0.04 0.027 0.122 0.045 ;
  END
END BUFx4_ASAP7_6t_SL

MACRO BUFx4q_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx4q_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.124 0.117 ;
        RECT 0.018 0.171 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.171 0.412 0.189 ;
        RECT 0.394 0.027 0.412 0.189 ;
        RECT 0.202 0.027 0.412 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.099 0.171 0.177 0.189 ;
      RECT 0.159 0.027 0.177 0.189 ;
      RECT 0.159 0.099 0.365 0.117 ;
      RECT 0.099 0.027 0.177 0.045 ;
  END
END BUFx4q_ASAP7_6t_SL

MACRO BUFx5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx5_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.011 0.099 0.078 0.117 ;
        RECT 0.011 0.135 0.066 0.153 ;
        RECT 0.011 0.063 0.066 0.081 ;
        RECT 0.011 0.063 0.029 0.153 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.171 0.414 0.189 ;
        RECT 0.396 0.027 0.414 0.189 ;
        RECT 0.148 0.027 0.414 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.171 0.122 0.189 ;
      RECT 0.104 0.027 0.122 0.189 ;
      RECT 0.104 0.099 0.365 0.117 ;
      RECT 0.04 0.027 0.122 0.045 ;
  END
END BUFx5_ASAP7_6t_SL

MACRO BUFx6q_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx6q_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.084 0.117 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.171 0.522 0.189 ;
        RECT 0.504 0.027 0.522 0.189 ;
        RECT 0.202 0.027 0.522 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.171 0.144 0.189 ;
      RECT 0.126 0.027 0.144 0.189 ;
      RECT 0.126 0.099 0.473 0.117 ;
      RECT 0.094 0.027 0.144 0.045 ;
  END
END BUFx6q_ASAP7_6t_SL

MACRO BUFx8_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx8_ASAP7_6t_SL 0 0 ;
  SIZE 0.648 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.095 0.117 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.648 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.171 0.63 0.189 ;
        RECT 0.612 0.027 0.63 0.189 ;
        RECT 0.202 0.027 0.63 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.171 0.144 0.189 ;
      RECT 0.126 0.027 0.144 0.189 ;
      RECT 0.126 0.099 0.581 0.117 ;
      RECT 0.094 0.027 0.144 0.045 ;
  END
END BUFx8_ASAP7_6t_SL

MACRO CKINVDCx10_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKINVDCx10_ASAP7_6t_SL 0 0 ;
  SIZE 1.296 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.071 0.099 1.17 0.117 ;
        RECT 1.12 0.027 1.138 0.117 ;
        RECT 0.018 0.027 1.138 0.045 ;
        RECT 0.747 0.099 0.814 0.117 ;
        RECT 0.796 0.027 0.814 0.117 ;
        RECT 0.374 0.099 0.441 0.117 ;
        RECT 0.374 0.027 0.392 0.117 ;
        RECT 0.018 0.099 0.117 0.117 ;
        RECT 0.018 0.171 0.068 0.189 ;
        RECT 0.018 0.027 0.037 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.296 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.296 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.171 1.224 0.189 ;
        RECT 1.206 0.027 1.224 0.189 ;
        RECT 1.174 0.027 1.224 0.045 ;
        RECT 1.028 0.063 1.094 0.081 ;
        RECT 1.028 0.063 1.046 0.189 ;
        RECT 0.704 0.063 0.77 0.081 ;
        RECT 0.704 0.063 0.722 0.189 ;
        RECT 0.466 0.063 0.484 0.189 ;
        RECT 0.418 0.063 0.484 0.081 ;
        RECT 0.142 0.063 0.16 0.189 ;
        RECT 0.094 0.063 0.16 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.936 0.099 0.992 0.117 ;
      RECT 0.936 0.063 0.954 0.117 ;
      RECT 0.85 0.063 1.002 0.081 ;
      RECT 0.831 0.135 0.986 0.153 ;
      RECT 0.882 0.099 0.9 0.153 ;
      RECT 0.842 0.099 0.9 0.117 ;
      RECT 0.526 0.135 0.675 0.153 ;
      RECT 0.612 0.099 0.63 0.153 ;
      RECT 0.612 0.099 0.67 0.117 ;
      RECT 0.52 0.099 0.576 0.117 ;
      RECT 0.558 0.063 0.576 0.117 ;
      RECT 0.51 0.063 0.662 0.081 ;
      RECT 0.202 0.135 0.357 0.153 ;
      RECT 0.288 0.099 0.306 0.153 ;
      RECT 0.288 0.099 0.346 0.117 ;
      RECT 0.196 0.099 0.252 0.117 ;
      RECT 0.234 0.063 0.252 0.117 ;
      RECT 0.186 0.063 0.338 0.081 ;
  END
END CKINVDCx10_ASAP7_6t_SL

MACRO CKINVDCx11_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKINVDCx11_ASAP7_6t_SL 0 0 ;
  SIZE 1.404 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.287 0.099 1.364 0.117 ;
        RECT 1.336 0.027 1.364 0.117 ;
        RECT 0.04 0.027 1.364 0.045 ;
        RECT 0.855 0.099 0.981 0.117 ;
        RECT 0.909 0.027 0.927 0.117 ;
        RECT 0.423 0.099 0.549 0.117 ;
        RECT 0.476 0.027 0.494 0.117 ;
        RECT 0.04 0.099 0.117 0.117 ;
        RECT 0.04 0.027 0.067 0.117 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.404 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.404 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.092 0.171 1.31 0.189 ;
        RECT 1.244 0.063 1.305 0.081 ;
        RECT 1.244 0.063 1.262 0.189 ;
        RECT 1.006 0.063 1.024 0.189 ;
        RECT 0.956 0.063 1.024 0.081 ;
        RECT 0.808 0.063 0.873 0.081 ;
        RECT 0.808 0.063 0.83 0.189 ;
        RECT 0.575 0.063 0.593 0.189 ;
        RECT 0.524 0.063 0.593 0.081 ;
        RECT 0.38 0.063 0.441 0.081 ;
        RECT 0.38 0.063 0.398 0.189 ;
        RECT 0.142 0.063 0.16 0.189 ;
        RECT 0.092 0.063 0.16 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.152 0.099 1.208 0.117 ;
      RECT 1.152 0.063 1.17 0.117 ;
      RECT 1.066 0.063 1.218 0.081 ;
      RECT 1.054 0.135 1.202 0.153 ;
      RECT 1.098 0.099 1.116 0.153 ;
      RECT 1.058 0.099 1.116 0.117 ;
      RECT 0.634 0.135 0.782 0.153 ;
      RECT 0.72 0.099 0.738 0.153 ;
      RECT 0.72 0.099 0.778 0.117 ;
      RECT 0.628 0.099 0.684 0.117 ;
      RECT 0.666 0.063 0.684 0.117 ;
      RECT 0.618 0.063 0.77 0.081 ;
      RECT 0.202 0.135 0.349 0.153 ;
      RECT 0.288 0.099 0.306 0.153 ;
      RECT 0.288 0.099 0.346 0.117 ;
      RECT 0.196 0.099 0.252 0.117 ;
      RECT 0.234 0.063 0.252 0.117 ;
      RECT 0.186 0.063 0.338 0.081 ;
  END
END CKINVDCx11_ASAP7_6t_SL

MACRO CKINVDCx12_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKINVDCx12_ASAP7_6t_SL 0 0 ;
  SIZE 1.404 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.281 0.099 1.354 0.117 ;
        RECT 1.336 0.027 1.354 0.117 ;
        RECT 0.049 0.027 1.354 0.045 ;
        RECT 0.85 0.099 0.986 0.117 ;
        RECT 0.909 0.027 0.927 0.117 ;
        RECT 0.418 0.099 0.554 0.117 ;
        RECT 0.476 0.027 0.494 0.117 ;
        RECT 0.049 0.099 0.122 0.117 ;
        RECT 0.049 0.027 0.067 0.117 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.404 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.404 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.092 0.171 1.311 0.189 ;
        RECT 1.237 0.063 1.31 0.081 ;
        RECT 1.237 0.063 1.255 0.189 ;
        RECT 1.011 0.063 1.029 0.189 ;
        RECT 0.956 0.063 1.029 0.081 ;
        RECT 0.803 0.063 0.878 0.081 ;
        RECT 0.803 0.063 0.823 0.189 ;
        RECT 0.583 0.063 0.603 0.189 ;
        RECT 0.524 0.063 0.603 0.081 ;
        RECT 0.372 0.063 0.446 0.081 ;
        RECT 0.372 0.063 0.39 0.189 ;
        RECT 0.152 0.063 0.17 0.189 ;
        RECT 0.092 0.063 0.17 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.152 0.099 1.209 0.117 ;
      RECT 1.152 0.063 1.17 0.117 ;
      RECT 1.059 0.063 1.21 0.081 ;
      RECT 1.059 0.135 1.202 0.153 ;
      RECT 1.098 0.099 1.116 0.153 ;
      RECT 1.059 0.099 1.116 0.117 ;
      RECT 0.634 0.135 0.775 0.153 ;
      RECT 0.72 0.099 0.738 0.153 ;
      RECT 0.72 0.099 0.775 0.117 ;
      RECT 0.628 0.099 0.684 0.117 ;
      RECT 0.666 0.063 0.684 0.117 ;
      RECT 0.628 0.063 0.77 0.081 ;
      RECT 0.202 0.135 0.346 0.153 ;
      RECT 0.288 0.099 0.306 0.153 ;
      RECT 0.288 0.099 0.346 0.117 ;
      RECT 0.196 0.099 0.252 0.117 ;
      RECT 0.234 0.063 0.252 0.117 ;
      RECT 0.196 0.063 0.338 0.081 ;
  END
END CKINVDCx12_ASAP7_6t_SL

MACRO CKINVDCx14_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKINVDCx14_ASAP7_6t_SL 0 0 ;
  SIZE 1.512 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.304 0.099 1.397 0.117 ;
        RECT 1.341 0.027 1.359 0.117 ;
        RECT 0.04 0.027 1.359 0.045 ;
        RECT 0.872 0.099 0.964 0.117 ;
        RECT 0.909 0.027 0.927 0.117 ;
        RECT 0.439 0.099 0.531 0.117 ;
        RECT 0.476 0.027 0.494 0.117 ;
        RECT 0.04 0.099 0.101 0.117 ;
        RECT 0.04 0.027 0.064 0.117 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.512 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.512 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 1.472 0.189 ;
        RECT 1.454 0.027 1.472 0.189 ;
        RECT 1.384 0.027 1.472 0.045 ;
        RECT 1.26 0.063 1.315 0.081 ;
        RECT 1.26 0.063 1.278 0.189 ;
        RECT 0.99 0.063 1.008 0.189 ;
        RECT 0.952 0.063 1.008 0.081 ;
        RECT 0.828 0.063 0.883 0.081 ;
        RECT 0.828 0.063 0.846 0.189 ;
        RECT 0.558 0.063 0.576 0.189 ;
        RECT 0.521 0.063 0.576 0.081 ;
        RECT 0.396 0.063 0.451 0.081 ;
        RECT 0.396 0.063 0.414 0.189 ;
        RECT 0.126 0.063 0.144 0.189 ;
        RECT 0.089 0.063 0.144 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.152 0.099 1.208 0.117 ;
      RECT 1.152 0.063 1.17 0.117 ;
      RECT 1.066 0.063 1.218 0.081 ;
      RECT 1.047 0.135 1.202 0.153 ;
      RECT 1.098 0.099 1.116 0.153 ;
      RECT 1.058 0.099 1.116 0.117 ;
      RECT 0.634 0.135 0.789 0.153 ;
      RECT 0.72 0.099 0.738 0.153 ;
      RECT 0.72 0.099 0.778 0.117 ;
      RECT 0.628 0.099 0.684 0.117 ;
      RECT 0.666 0.063 0.684 0.117 ;
      RECT 0.618 0.063 0.77 0.081 ;
      RECT 0.202 0.135 0.357 0.153 ;
      RECT 0.288 0.099 0.306 0.153 ;
      RECT 0.288 0.099 0.346 0.117 ;
      RECT 0.196 0.099 0.252 0.117 ;
      RECT 0.234 0.063 0.252 0.117 ;
      RECT 0.186 0.063 0.338 0.081 ;
  END
END CKINVDCx14_ASAP7_6t_SL

MACRO CKINVDCx16_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKINVDCx16_ASAP7_6t_SL 0 0 ;
  SIZE 1.62 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.552 0.171 1.602 0.189 ;
        RECT 1.584 0.027 1.602 0.189 ;
        RECT 1.423 0.099 1.602 0.117 ;
        RECT 0.152 0.027 1.602 0.045 ;
        RECT 0.98 0.099 1.072 0.117 ;
        RECT 1.017 0.027 1.035 0.117 ;
        RECT 0.547 0.099 0.639 0.117 ;
        RECT 0.584 0.027 0.602 0.117 ;
        RECT 0.118 0.099 0.207 0.117 ;
        RECT 0.152 0.027 0.17 0.117 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.62 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.62 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.057 0.171 1.521 0.189 ;
        RECT 1.368 0.063 1.521 0.081 ;
        RECT 1.368 0.063 1.386 0.189 ;
        RECT 1.098 0.063 1.116 0.189 ;
        RECT 1.061 0.063 1.116 0.081 ;
        RECT 0.936 0.063 0.991 0.081 ;
        RECT 0.936 0.063 0.954 0.189 ;
        RECT 0.666 0.063 0.684 0.189 ;
        RECT 0.628 0.063 0.684 0.081 ;
        RECT 0.504 0.063 0.559 0.081 ;
        RECT 0.504 0.063 0.522 0.189 ;
        RECT 0.234 0.063 0.252 0.189 ;
        RECT 0.196 0.063 0.252 0.081 ;
        RECT 0.057 0.027 0.122 0.045 ;
        RECT 0.057 0.027 0.075 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.26 0.099 1.316 0.117 ;
      RECT 1.26 0.063 1.278 0.117 ;
      RECT 1.174 0.063 1.326 0.081 ;
      RECT 1.155 0.135 1.31 0.153 ;
      RECT 1.206 0.099 1.224 0.153 ;
      RECT 1.166 0.099 1.224 0.117 ;
      RECT 0.742 0.135 0.897 0.153 ;
      RECT 0.828 0.099 0.846 0.153 ;
      RECT 0.828 0.099 0.886 0.117 ;
      RECT 0.736 0.099 0.792 0.117 ;
      RECT 0.774 0.063 0.792 0.117 ;
      RECT 0.726 0.063 0.878 0.081 ;
      RECT 0.31 0.135 0.465 0.153 ;
      RECT 0.396 0.099 0.414 0.153 ;
      RECT 0.396 0.099 0.454 0.117 ;
      RECT 0.304 0.099 0.36 0.117 ;
      RECT 0.342 0.063 0.36 0.117 ;
      RECT 0.294 0.063 0.446 0.081 ;
  END
END CKINVDCx16_ASAP7_6t_SL

MACRO CKINVDCx20_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKINVDCx20_ASAP7_6t_SL 0 0 ;
  SIZE 2.052 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.843 0.099 1.937 0.117 ;
        RECT 1.88 0.027 1.904 0.117 ;
        RECT 0.148 0.027 1.904 0.045 ;
        RECT 1.412 0.099 1.505 0.117 ;
        RECT 1.449 0.027 1.467 0.117 ;
        RECT 0.98 0.099 1.072 0.117 ;
        RECT 1.017 0.027 1.035 0.117 ;
        RECT 0.547 0.099 0.64 0.117 ;
        RECT 0.585 0.027 0.603 0.117 ;
        RECT 0.126 0.099 0.208 0.117 ;
        RECT 0.148 0.027 0.171 0.117 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 2.052 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 2.052 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.04 0.171 2.012 0.189 ;
        RECT 1.994 0.027 2.012 0.189 ;
        RECT 1.93 0.027 2.012 0.045 ;
        RECT 1.8 0.063 1.855 0.081 ;
        RECT 1.8 0.063 1.818 0.189 ;
        RECT 1.53 0.063 1.548 0.189 ;
        RECT 1.493 0.063 1.548 0.081 ;
        RECT 1.368 0.063 1.423 0.081 ;
        RECT 1.368 0.063 1.386 0.189 ;
        RECT 1.098 0.063 1.116 0.189 ;
        RECT 1.061 0.063 1.116 0.081 ;
        RECT 0.936 0.063 0.991 0.081 ;
        RECT 0.936 0.063 0.954 0.189 ;
        RECT 0.666 0.063 0.684 0.189 ;
        RECT 0.629 0.063 0.684 0.081 ;
        RECT 0.504 0.063 0.559 0.081 ;
        RECT 0.504 0.063 0.522 0.189 ;
        RECT 0.234 0.063 0.252 0.189 ;
        RECT 0.197 0.063 0.252 0.081 ;
        RECT 0.04 0.027 0.122 0.045 ;
        RECT 0.04 0.027 0.058 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.692 0.099 1.748 0.117 ;
      RECT 1.692 0.063 1.71 0.117 ;
      RECT 1.606 0.063 1.758 0.081 ;
      RECT 1.587 0.135 1.742 0.153 ;
      RECT 1.638 0.099 1.656 0.153 ;
      RECT 1.598 0.099 1.656 0.117 ;
      RECT 1.26 0.099 1.316 0.117 ;
      RECT 1.26 0.063 1.278 0.117 ;
      RECT 1.174 0.063 1.326 0.081 ;
      RECT 1.155 0.135 1.31 0.153 ;
      RECT 1.206 0.099 1.224 0.153 ;
      RECT 1.166 0.099 1.224 0.117 ;
      RECT 0.742 0.135 0.897 0.153 ;
      RECT 0.828 0.099 0.846 0.153 ;
      RECT 0.828 0.099 0.886 0.117 ;
      RECT 0.736 0.099 0.792 0.117 ;
      RECT 0.774 0.063 0.792 0.117 ;
      RECT 0.726 0.063 0.878 0.081 ;
      RECT 0.31 0.135 0.465 0.153 ;
      RECT 0.396 0.099 0.414 0.153 ;
      RECT 0.396 0.099 0.454 0.117 ;
      RECT 0.304 0.099 0.36 0.117 ;
      RECT 0.342 0.063 0.36 0.117 ;
      RECT 0.294 0.063 0.446 0.081 ;
  END
END CKINVDCx20_ASAP7_6t_SL

MACRO CKINVDCx5p5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKINVDCx5p5_ASAP7_6t_SL 0 0 ;
  SIZE 1.134 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.099 1.084 0.117 ;
        RECT 1.066 0.027 1.084 0.117 ;
        RECT 0.094 0.027 1.084 0.045 ;
        RECT 0.688 0.099 0.76 0.117 ;
        RECT 0.742 0.027 0.76 0.117 ;
        RECT 0.32 0.099 0.392 0.117 ;
        RECT 0.32 0.027 0.338 0.117 ;
        RECT 0.067 0.099 0.112 0.117 ;
        RECT 0.094 0.027 0.112 0.117 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.134 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.134 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.023 0.171 1.04 0.189 ;
        RECT 0.969 0.063 1.04 0.081 ;
        RECT 0.969 0.063 0.987 0.189 ;
        RECT 0.645 0.063 0.716 0.081 ;
        RECT 0.645 0.063 0.663 0.189 ;
        RECT 0.417 0.063 0.435 0.189 ;
        RECT 0.364 0.063 0.435 0.081 ;
        RECT 0.023 0.027 0.068 0.045 ;
        RECT 0.023 0.027 0.042 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.882 0.099 0.938 0.117 ;
      RECT 0.882 0.063 0.9 0.117 ;
      RECT 0.796 0.063 0.944 0.081 ;
      RECT 0.777 0.135 0.932 0.153 ;
      RECT 0.828 0.099 0.846 0.153 ;
      RECT 0.788 0.099 0.846 0.117 ;
      RECT 0.472 0.135 0.616 0.153 ;
      RECT 0.558 0.099 0.576 0.153 ;
      RECT 0.558 0.099 0.616 0.117 ;
      RECT 0.466 0.099 0.522 0.117 ;
      RECT 0.504 0.063 0.522 0.117 ;
      RECT 0.463 0.063 0.608 0.081 ;
      RECT 0.148 0.135 0.303 0.153 ;
      RECT 0.234 0.099 0.252 0.153 ;
      RECT 0.234 0.099 0.292 0.117 ;
      RECT 0.142 0.099 0.198 0.117 ;
      RECT 0.18 0.063 0.198 0.117 ;
      RECT 0.142 0.063 0.284 0.081 ;
  END
END CKINVDCx5p5_ASAP7_6t_SL

MACRO CKINVDCx6p5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKINVDCx6p5_ASAP7_6t_SL 0 0 ;
  SIZE 1.242 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.071 0.099 1.163 0.117 ;
        RECT 0.04 0.027 1.148 0.045 ;
        RECT 1.12 0.027 1.138 0.117 ;
        RECT 0.747 0.099 0.814 0.117 ;
        RECT 0.796 0.027 0.814 0.117 ;
        RECT 0.374 0.099 0.441 0.117 ;
        RECT 0.374 0.027 0.392 0.117 ;
        RECT 0.04 0.099 0.117 0.117 ;
        RECT 0.04 0.027 0.068 0.117 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.242 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.242 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 1.216 0.189 ;
        RECT 1.198 0.063 1.216 0.189 ;
        RECT 1.174 0.063 1.216 0.081 ;
        RECT 1.028 0.063 1.094 0.081 ;
        RECT 1.028 0.063 1.046 0.189 ;
        RECT 0.702 0.063 0.77 0.081 ;
        RECT 0.702 0.063 0.72 0.189 ;
        RECT 0.467 0.063 0.485 0.189 ;
        RECT 0.418 0.063 0.485 0.081 ;
        RECT 0.144 0.063 0.162 0.189 ;
        RECT 0.094 0.063 0.162 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.936 0.099 0.992 0.117 ;
      RECT 0.936 0.063 0.954 0.117 ;
      RECT 0.85 0.063 1.002 0.081 ;
      RECT 0.831 0.135 0.986 0.153 ;
      RECT 0.882 0.099 0.9 0.153 ;
      RECT 0.842 0.099 0.9 0.117 ;
      RECT 0.526 0.135 0.676 0.153 ;
      RECT 0.612 0.099 0.63 0.153 ;
      RECT 0.612 0.099 0.67 0.117 ;
      RECT 0.52 0.099 0.576 0.117 ;
      RECT 0.558 0.063 0.576 0.117 ;
      RECT 0.511 0.063 0.662 0.081 ;
      RECT 0.202 0.135 0.357 0.153 ;
      RECT 0.288 0.099 0.306 0.153 ;
      RECT 0.288 0.099 0.346 0.117 ;
      RECT 0.196 0.099 0.252 0.117 ;
      RECT 0.234 0.063 0.252 0.117 ;
      RECT 0.189 0.063 0.338 0.081 ;
  END
END CKINVDCx6p5_ASAP7_6t_SL

MACRO CKINVDCx8_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKINVDCx8_ASAP7_6t_SL 0 0 ;
  SIZE 1.188 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.018 0.099 1.09 0.117 ;
        RECT 1.018 0.027 1.036 0.117 ;
        RECT 0.027 0.027 1.036 0.045 ;
        RECT 0.747 0.099 0.817 0.117 ;
        RECT 0.799 0.027 0.817 0.117 ;
        RECT 0.371 0.099 0.441 0.117 ;
        RECT 0.371 0.027 0.389 0.117 ;
        RECT 0.027 0.099 0.085 0.117 ;
        RECT 0.027 0.171 0.068 0.189 ;
        RECT 0.027 0.027 0.045 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.188 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.188 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.171 1.137 0.189 ;
        RECT 1.119 0.027 1.137 0.189 ;
        RECT 1.066 0.027 1.137 0.045 ;
        RECT 0.704 0.063 0.771 0.081 ;
        RECT 0.704 0.063 0.722 0.189 ;
        RECT 0.466 0.063 0.484 0.189 ;
        RECT 0.417 0.063 0.484 0.081 ;
        RECT 0.126 0.063 0.144 0.189 ;
        RECT 0.094 0.063 0.144 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.936 0.099 0.992 0.117 ;
      RECT 0.936 0.063 0.954 0.117 ;
      RECT 0.85 0.063 0.993 0.081 ;
      RECT 0.84 0.135 0.986 0.153 ;
      RECT 0.882 0.099 0.9 0.153 ;
      RECT 0.842 0.099 0.9 0.117 ;
      RECT 0.526 0.135 0.679 0.153 ;
      RECT 0.612 0.099 0.63 0.153 ;
      RECT 0.612 0.099 0.67 0.117 ;
      RECT 0.52 0.099 0.576 0.117 ;
      RECT 0.558 0.063 0.576 0.117 ;
      RECT 0.51 0.063 0.662 0.081 ;
      RECT 0.202 0.135 0.352 0.153 ;
      RECT 0.288 0.099 0.306 0.153 ;
      RECT 0.288 0.099 0.346 0.117 ;
      RECT 0.196 0.099 0.252 0.117 ;
      RECT 0.234 0.063 0.252 0.117 ;
      RECT 0.186 0.063 0.338 0.081 ;
  END
END CKINVDCx8_ASAP7_6t_SL

MACRO CKINVDCx9p5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CKINVDCx9p5_ASAP7_6t_SL 0 0 ;
  SIZE 1.512 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.287 0.099 1.413 0.117 ;
        RECT 1.339 0.027 1.364 0.117 ;
        RECT 0.04 0.027 1.364 0.045 ;
        RECT 0.855 0.099 0.981 0.117 ;
        RECT 0.909 0.027 0.927 0.117 ;
        RECT 0.423 0.099 0.549 0.117 ;
        RECT 0.476 0.027 0.494 0.117 ;
        RECT 0.04 0.099 0.117 0.117 ;
        RECT 0.04 0.027 0.064 0.117 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.512 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.512 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.04 0.171 1.472 0.189 ;
        RECT 1.454 0.063 1.472 0.189 ;
        RECT 1.39 0.063 1.472 0.081 ;
        RECT 1.244 0.063 1.31 0.081 ;
        RECT 1.244 0.063 1.262 0.189 ;
        RECT 1.006 0.063 1.024 0.189 ;
        RECT 0.958 0.063 1.024 0.081 ;
        RECT 0.812 0.063 0.878 0.081 ;
        RECT 0.812 0.063 0.83 0.189 ;
        RECT 0.574 0.063 0.592 0.189 ;
        RECT 0.526 0.063 0.592 0.081 ;
        RECT 0.38 0.063 0.446 0.081 ;
        RECT 0.38 0.063 0.398 0.189 ;
        RECT 0.142 0.063 0.16 0.189 ;
        RECT 0.089 0.063 0.16 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.152 0.099 1.208 0.117 ;
      RECT 1.152 0.063 1.17 0.117 ;
      RECT 1.066 0.063 1.218 0.081 ;
      RECT 1.055 0.135 1.202 0.153 ;
      RECT 1.098 0.099 1.116 0.153 ;
      RECT 1.058 0.099 1.116 0.117 ;
      RECT 0.634 0.135 0.78 0.153 ;
      RECT 0.72 0.099 0.738 0.153 ;
      RECT 0.72 0.099 0.778 0.117 ;
      RECT 0.628 0.099 0.684 0.117 ;
      RECT 0.666 0.063 0.684 0.117 ;
      RECT 0.618 0.063 0.77 0.081 ;
      RECT 0.202 0.135 0.348 0.153 ;
      RECT 0.288 0.099 0.306 0.153 ;
      RECT 0.288 0.099 0.346 0.117 ;
      RECT 0.196 0.099 0.252 0.117 ;
      RECT 0.234 0.063 0.252 0.117 ;
      RECT 0.186 0.063 0.338 0.081 ;
  END
END CKINVDCx9p5_ASAP7_6t_SL

MACRO DECAPx10_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DECAPx10_ASAP7_6t_SL 0 0 ;
  SIZE 1.188 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.188 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.188 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.558 0.045 0.576 0.117 ;
      RECT 0.558 0.045 1.148 0.063 ;
      RECT 0.04 0.153 0.63 0.171 ;
      RECT 0.612 0.099 0.63 0.171 ;
  END
END DECAPx10_ASAP7_6t_SL

MACRO DECAPx1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DECAPx1_ASAP7_6t_SL 0 0 ;
  SIZE 0.216 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.216 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.216 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.094 0.153 0.144 0.171 ;
      RECT 0.126 0.099 0.144 0.171 ;
      RECT 0.072 0.045 0.09 0.117 ;
      RECT 0.072 0.045 0.117 0.063 ;
  END
END DECAPx1_ASAP7_6t_SL

MACRO DECAPx2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DECAPx2_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.126 0.045 0.144 0.117 ;
      RECT 0.126 0.045 0.284 0.063 ;
      RECT 0.04 0.153 0.198 0.171 ;
      RECT 0.18 0.099 0.198 0.171 ;
  END
END DECAPx2_ASAP7_6t_SL

MACRO DECAPx2b_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DECAPx2b_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.094 0.135 0.249 0.153 ;
      RECT 0.18 0.099 0.198 0.153 ;
      RECT 0.18 0.099 0.238 0.117 ;
      RECT 0.088 0.099 0.144 0.117 ;
      RECT 0.126 0.063 0.144 0.117 ;
      RECT 0.078 0.063 0.23 0.081 ;
  END
END DECAPx2b_ASAP7_6t_SL

MACRO DECAPx4_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DECAPx4_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.234 0.045 0.252 0.117 ;
      RECT 0.234 0.045 0.5 0.063 ;
      RECT 0.04 0.153 0.306 0.171 ;
      RECT 0.288 0.099 0.306 0.171 ;
  END
END DECAPx4_ASAP7_6t_SL

MACRO DECAPx6_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DECAPx6_ASAP7_6t_SL 0 0 ;
  SIZE 0.756 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.756 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.756 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.342 0.045 0.36 0.117 ;
      RECT 0.342 0.045 0.716 0.063 ;
      RECT 0.04 0.153 0.414 0.171 ;
      RECT 0.396 0.099 0.414 0.171 ;
  END
END DECAPx6_ASAP7_6t_SL

MACRO DFFARHQNx1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFARHQNx1_ASAP7_6t_SL 0 0 ;
  SIZE 1.296 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.052 0.171 0.135 0.189 ;
        RECT 0.052 0.027 0.135 0.045 ;
        RECT 0.052 0.099 0.09 0.117 ;
        RECT 0.052 0.027 0.07 0.189 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.27 0.027 0.345 0.045 ;
        RECT 0.191 0.171 0.309 0.189 ;
        RECT 0.27 0.099 0.306 0.117 ;
        RECT 0.27 0.027 0.288 0.189 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.213 0.171 1.278 0.189 ;
        RECT 1.26 0.027 1.278 0.189 ;
        RECT 1.213 0.027 1.278 0.045 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.296 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.296 0.009 ;
    END
  END VSS
  PIN RESETN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.526 0.027 1.148 0.045 ;
      LAYER M1 ;
        RECT 1.111 0.027 1.152 0.045 ;
        RECT 1.111 0.027 1.129 0.098 ;
        RECT 0.505 0.027 0.561 0.045 ;
        RECT 0.505 0.027 0.523 0.088 ;
      LAYER V1 ;
        RECT 0.531 0.027 0.549 0.045 ;
        RECT 1.125 0.027 1.143 0.045 ;
    END
  END RESETN
  OBS
    LAYER M1 ;
      RECT 1.206 0.063 1.224 0.125 ;
      RECT 1.192 0.063 1.229 0.081 ;
      RECT 1.069 0.171 1.149 0.189 ;
      RECT 1.069 0.027 1.087 0.189 ;
      RECT 0.936 0.027 0.954 0.088 ;
      RECT 0.936 0.027 1.087 0.045 ;
      RECT 0.954 0.135 0.988 0.153 ;
      RECT 0.954 0.113 0.974 0.153 ;
      RECT 0.907 0.113 0.974 0.131 ;
      RECT 0.855 0.13 0.873 0.175 ;
      RECT 0.864 0.027 0.882 0.151 ;
      RECT 0.864 0.063 0.904 0.081 ;
      RECT 0.796 0.027 0.882 0.045 ;
      RECT 0.828 0.063 0.846 0.104 ;
      RECT 0.808 0.063 0.846 0.081 ;
      RECT 0.749 0.171 0.824 0.189 ;
      RECT 0.749 0.027 0.767 0.189 ;
      RECT 0.614 0.027 0.632 0.132 ;
      RECT 0.614 0.027 0.767 0.045 ;
      RECT 0.785 0.135 0.822 0.153 ;
      RECT 0.785 0.108 0.803 0.153 ;
      RECT 0.542 0.135 0.58 0.153 ;
      RECT 0.503 0.119 0.569 0.137 ;
      RECT 0.354 0.171 0.449 0.189 ;
      RECT 0.431 0.054 0.449 0.189 ;
      RECT 0.393 0.063 0.411 0.126 ;
      RECT 0.374 0.063 0.411 0.081 ;
      RECT 0.322 0.135 0.36 0.153 ;
      RECT 0.342 0.098 0.36 0.153 ;
      RECT 0.182 0.135 0.252 0.153 ;
      RECT 0.234 0.063 0.252 0.153 ;
      RECT 0.195 0.063 0.252 0.081 ;
      RECT 0.126 0.063 0.144 0.126 ;
      RECT 0.111 0.063 0.154 0.081 ;
      RECT 0.66 0.099 0.719 0.117 ;
      RECT 0.477 0.171 0.623 0.189 ;
      RECT 0.016 0.049 0.034 0.167 ;
    LAYER M2 ;
      RECT 0.882 0.063 1.229 0.081 ;
      RECT 0.202 0.135 0.986 0.153 ;
      RECT 0.016 0.063 0.839 0.081 ;
      RECT 0.426 0.099 0.704 0.117 ;
    LAYER V1 ;
      RECT 1.206 0.063 1.224 0.081 ;
      RECT 0.963 0.135 0.981 0.153 ;
      RECT 0.882 0.063 0.9 0.081 ;
      RECT 0.821 0.063 0.839 0.081 ;
      RECT 0.79 0.135 0.808 0.153 ;
      RECT 0.676 0.099 0.694 0.117 ;
      RECT 0.551 0.135 0.569 0.153 ;
      RECT 0.431 0.099 0.449 0.117 ;
      RECT 0.385 0.063 0.403 0.081 ;
      RECT 0.333 0.135 0.351 0.153 ;
      RECT 0.207 0.135 0.225 0.153 ;
      RECT 0.126 0.063 0.144 0.081 ;
      RECT 0.016 0.063 0.034 0.081 ;
  END
END DFFARHQNx1_ASAP7_6t_SL

MACRO DFFASHQNx1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFASHQNx1_ASAP7_6t_SL 0 0 ;
  SIZE 1.296 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.052 0.171 0.135 0.189 ;
        RECT 0.052 0.027 0.135 0.045 ;
        RECT 0.052 0.099 0.09 0.117 ;
        RECT 0.052 0.027 0.07 0.189 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.27 0.027 0.345 0.045 ;
        RECT 0.191 0.171 0.309 0.189 ;
        RECT 0.27 0.099 0.306 0.117 ;
        RECT 0.27 0.027 0.288 0.189 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.213 0.171 1.278 0.189 ;
        RECT 1.26 0.027 1.278 0.189 ;
        RECT 1.213 0.027 1.278 0.045 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.296 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.296 0.009 ;
    END
  END VSS
  PIN SETN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.708 0.099 1.092 0.117 ;
      LAYER M1 ;
        RECT 1.069 0.07 1.087 0.142 ;
        RECT 0.99 0.07 1.087 0.088 ;
        RECT 0.684 0.171 0.731 0.189 ;
        RECT 0.713 0.094 0.731 0.189 ;
      LAYER V1 ;
        RECT 0.713 0.099 0.731 0.117 ;
        RECT 1.069 0.099 1.087 0.117 ;
    END
  END SETN
  OBS
    LAYER M1 ;
      RECT 1.206 0.063 1.224 0.125 ;
      RECT 1.192 0.063 1.229 0.081 ;
      RECT 1.066 0.171 1.14 0.189 ;
      RECT 1.122 0.027 1.14 0.189 ;
      RECT 0.936 0.027 0.954 0.088 ;
      RECT 0.936 0.027 1.14 0.045 ;
      RECT 0.954 0.135 1.022 0.153 ;
      RECT 0.954 0.113 0.974 0.153 ;
      RECT 0.907 0.113 0.974 0.131 ;
      RECT 0.855 0.13 0.873 0.175 ;
      RECT 0.864 0.027 0.882 0.151 ;
      RECT 0.864 0.063 0.904 0.081 ;
      RECT 0.796 0.027 0.882 0.045 ;
      RECT 0.828 0.063 0.846 0.104 ;
      RECT 0.808 0.063 0.846 0.081 ;
      RECT 0.749 0.171 0.824 0.189 ;
      RECT 0.749 0.027 0.767 0.189 ;
      RECT 0.56 0.135 0.662 0.153 ;
      RECT 0.56 0.027 0.578 0.153 ;
      RECT 0.56 0.027 0.767 0.045 ;
      RECT 0.785 0.135 0.822 0.153 ;
      RECT 0.785 0.108 0.803 0.153 ;
      RECT 0.467 0.135 0.526 0.153 ;
      RECT 0.467 0.108 0.485 0.153 ;
      RECT 0.354 0.171 0.449 0.189 ;
      RECT 0.431 0.054 0.449 0.189 ;
      RECT 0.393 0.063 0.411 0.126 ;
      RECT 0.374 0.063 0.411 0.081 ;
      RECT 0.322 0.135 0.36 0.153 ;
      RECT 0.342 0.098 0.36 0.153 ;
      RECT 0.182 0.135 0.252 0.153 ;
      RECT 0.234 0.063 0.252 0.153 ;
      RECT 0.195 0.063 0.252 0.081 ;
      RECT 0.126 0.063 0.144 0.126 ;
      RECT 0.111 0.063 0.154 0.081 ;
      RECT 0.904 0.171 1.035 0.189 ;
      RECT 0.606 0.099 0.665 0.117 ;
      RECT 0.016 0.049 0.034 0.167 ;
    LAYER M2 ;
      RECT 0.882 0.063 1.231 0.081 ;
      RECT 0.202 0.135 1.013 0.153 ;
      RECT 0.016 0.063 0.839 0.081 ;
      RECT 0.426 0.099 0.65 0.117 ;
    LAYER V1 ;
      RECT 1.206 0.063 1.224 0.081 ;
      RECT 0.99 0.135 1.008 0.153 ;
      RECT 0.882 0.063 0.9 0.081 ;
      RECT 0.821 0.063 0.839 0.081 ;
      RECT 0.79 0.135 0.808 0.153 ;
      RECT 0.622 0.099 0.64 0.117 ;
      RECT 0.497 0.135 0.515 0.153 ;
      RECT 0.431 0.099 0.449 0.117 ;
      RECT 0.385 0.063 0.403 0.081 ;
      RECT 0.333 0.135 0.351 0.153 ;
      RECT 0.207 0.135 0.225 0.153 ;
      RECT 0.126 0.063 0.144 0.081 ;
      RECT 0.016 0.063 0.034 0.081 ;
  END
END DFFASHQNx1_ASAP7_6t_SL

MACRO DFFASRHQNx1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFASRHQNx1_ASAP7_6t_SL 0 0 ;
  SIZE 1.404 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.052 0.171 0.135 0.189 ;
        RECT 0.052 0.027 0.135 0.045 ;
        RECT 0.052 0.099 0.09 0.117 ;
        RECT 0.052 0.027 0.07 0.189 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.27 0.027 0.345 0.045 ;
        RECT 0.191 0.171 0.309 0.189 ;
        RECT 0.27 0.099 0.306 0.117 ;
        RECT 0.27 0.027 0.288 0.189 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.321 0.171 1.386 0.189 ;
        RECT 1.368 0.027 1.386 0.189 ;
        RECT 1.321 0.027 1.386 0.045 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.404 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.404 0.009 ;
    END
  END VSS
  PIN RESETN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.526 0.027 1.256 0.045 ;
      LAYER M1 ;
        RECT 1.219 0.027 1.26 0.045 ;
        RECT 1.219 0.027 1.237 0.098 ;
        RECT 0.505 0.027 0.561 0.045 ;
        RECT 0.505 0.027 0.523 0.088 ;
      LAYER V1 ;
        RECT 0.531 0.027 0.549 0.045 ;
        RECT 1.233 0.027 1.251 0.045 ;
    END
  END RESETN
  PIN SETN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.762 0.099 1.164 0.117 ;
      LAYER M1 ;
        RECT 1.141 0.07 1.159 0.142 ;
        RECT 1.044 0.07 1.159 0.088 ;
        RECT 0.738 0.171 0.785 0.189 ;
        RECT 0.767 0.094 0.785 0.189 ;
      LAYER V1 ;
        RECT 0.767 0.099 0.785 0.117 ;
        RECT 1.141 0.099 1.159 0.117 ;
    END
  END SETN
  OBS
    LAYER M1 ;
      RECT 1.314 0.063 1.332 0.125 ;
      RECT 1.3 0.063 1.337 0.081 ;
      RECT 1.177 0.171 1.257 0.189 ;
      RECT 1.177 0.027 1.195 0.189 ;
      RECT 0.99 0.027 1.008 0.088 ;
      RECT 0.99 0.027 1.195 0.045 ;
      RECT 1.008 0.135 1.076 0.153 ;
      RECT 1.008 0.113 1.028 0.153 ;
      RECT 0.961 0.113 1.028 0.131 ;
      RECT 0.909 0.13 0.927 0.175 ;
      RECT 0.918 0.027 0.936 0.151 ;
      RECT 0.918 0.063 0.958 0.081 ;
      RECT 0.85 0.027 0.936 0.045 ;
      RECT 0.882 0.063 0.9 0.104 ;
      RECT 0.862 0.063 0.9 0.081 ;
      RECT 0.803 0.171 0.878 0.189 ;
      RECT 0.803 0.027 0.821 0.189 ;
      RECT 0.614 0.135 0.716 0.153 ;
      RECT 0.614 0.027 0.632 0.153 ;
      RECT 0.614 0.027 0.821 0.045 ;
      RECT 0.839 0.135 0.876 0.153 ;
      RECT 0.839 0.108 0.857 0.153 ;
      RECT 0.542 0.135 0.58 0.153 ;
      RECT 0.503 0.119 0.569 0.137 ;
      RECT 0.354 0.171 0.449 0.189 ;
      RECT 0.431 0.054 0.449 0.189 ;
      RECT 0.393 0.063 0.411 0.126 ;
      RECT 0.374 0.063 0.411 0.081 ;
      RECT 0.322 0.135 0.36 0.153 ;
      RECT 0.342 0.098 0.36 0.153 ;
      RECT 0.182 0.135 0.252 0.153 ;
      RECT 0.234 0.063 0.252 0.153 ;
      RECT 0.195 0.063 0.252 0.081 ;
      RECT 0.126 0.063 0.144 0.126 ;
      RECT 0.111 0.063 0.154 0.081 ;
      RECT 0.958 0.171 1.094 0.189 ;
      RECT 0.66 0.099 0.719 0.117 ;
      RECT 0.477 0.171 0.623 0.189 ;
      RECT 0.016 0.049 0.034 0.167 ;
    LAYER M2 ;
      RECT 0.936 0.063 1.337 0.081 ;
      RECT 0.202 0.135 1.067 0.153 ;
      RECT 0.016 0.063 0.893 0.081 ;
      RECT 0.426 0.099 0.704 0.117 ;
    LAYER V1 ;
      RECT 1.314 0.063 1.332 0.081 ;
      RECT 1.044 0.135 1.062 0.153 ;
      RECT 0.936 0.063 0.954 0.081 ;
      RECT 0.875 0.063 0.893 0.081 ;
      RECT 0.844 0.135 0.862 0.153 ;
      RECT 0.676 0.099 0.694 0.117 ;
      RECT 0.551 0.135 0.569 0.153 ;
      RECT 0.431 0.099 0.449 0.117 ;
      RECT 0.385 0.063 0.403 0.081 ;
      RECT 0.333 0.135 0.351 0.153 ;
      RECT 0.207 0.135 0.225 0.153 ;
      RECT 0.126 0.063 0.144 0.081 ;
      RECT 0.016 0.063 0.034 0.081 ;
  END
END DFFASRHQNx1_ASAP7_6t_SL

MACRO DFFHQNx1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNx1_ASAP7_6t_SL 0 0 ;
  SIZE 1.08 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.176 0.189 ;
        RECT 0.094 0.027 0.176 0.045 ;
        RECT 0.094 0.128 0.117 0.189 ;
        RECT 0.072 0.065 0.115 0.083 ;
        RECT 0.094 0.027 0.115 0.083 ;
        RECT 0.072 0.128 0.117 0.146 ;
        RECT 0.072 0.065 0.09 0.146 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.27 0.027 0.392 0.045 ;
        RECT 0.251 0.171 0.338 0.189 ;
        RECT 0.27 0.027 0.288 0.189 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.953 0.171 1.062 0.189 ;
        RECT 1.044 0.027 1.062 0.189 ;
        RECT 0.953 0.027 1.062 0.045 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.08 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.08 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.881 0.063 0.899 0.126 ;
      RECT 0.862 0.063 0.899 0.081 ;
      RECT 0.81 0.171 0.878 0.189 ;
      RECT 0.81 0.027 0.828 0.189 ;
      RECT 0.769 0.07 0.828 0.088 ;
      RECT 0.809 0.027 0.828 0.088 ;
      RECT 0.809 0.027 0.878 0.045 ;
      RECT 0.688 0.17 0.738 0.188 ;
      RECT 0.72 0.027 0.738 0.188 ;
      RECT 0.634 0.027 0.738 0.045 ;
      RECT 0.666 0.063 0.684 0.123 ;
      RECT 0.654 0.063 0.694 0.081 ;
      RECT 0.601 0.135 0.64 0.153 ;
      RECT 0.612 0.094 0.63 0.153 ;
      RECT 0.522 0.171 0.628 0.189 ;
      RECT 0.522 0.047 0.54 0.189 ;
      RECT 0.494 0.077 0.54 0.095 ;
      RECT 0.522 0.047 0.603 0.065 ;
      RECT 0.369 0.171 0.464 0.189 ;
      RECT 0.446 0.027 0.464 0.189 ;
      RECT 0.423 0.027 0.464 0.045 ;
      RECT 0.396 0.063 0.414 0.126 ;
      RECT 0.377 0.063 0.414 0.081 ;
      RECT 0.306 0.135 0.377 0.153 ;
      RECT 0.306 0.099 0.324 0.153 ;
      RECT 0.306 0.099 0.368 0.117 ;
      RECT 0.201 0.112 0.219 0.158 ;
      RECT 0.201 0.112 0.244 0.13 ;
      RECT 0.225 0.027 0.244 0.13 ;
      RECT 0.207 0.027 0.244 0.045 ;
      RECT 0.143 0.063 0.161 0.117 ;
      RECT 0.143 0.063 0.183 0.081 ;
      RECT 0.016 0.171 0.068 0.189 ;
      RECT 0.016 0.027 0.034 0.189 ;
      RECT 0.016 0.027 0.063 0.045 ;
      RECT 0.774 0.113 0.792 0.172 ;
      RECT 0.558 0.094 0.576 0.144 ;
      RECT 0.486 0.126 0.504 0.172 ;
    LAYER M2 ;
      RECT 0.72 0.063 0.899 0.081 ;
      RECT 0.196 0.135 0.797 0.153 ;
      RECT 0.016 0.063 0.684 0.081 ;
      RECT 0.446 0.099 0.576 0.117 ;
    LAYER V1 ;
      RECT 0.876 0.063 0.894 0.081 ;
      RECT 0.774 0.135 0.792 0.153 ;
      RECT 0.72 0.063 0.738 0.081 ;
      RECT 0.666 0.063 0.684 0.081 ;
      RECT 0.612 0.135 0.63 0.153 ;
      RECT 0.558 0.099 0.576 0.117 ;
      RECT 0.486 0.135 0.504 0.153 ;
      RECT 0.446 0.099 0.464 0.117 ;
      RECT 0.391 0.063 0.409 0.081 ;
      RECT 0.315 0.135 0.333 0.153 ;
      RECT 0.201 0.135 0.219 0.153 ;
      RECT 0.153 0.063 0.171 0.081 ;
      RECT 0.016 0.063 0.034 0.081 ;
  END
END DFFHQNx1_ASAP7_6t_SL

MACRO DFFHQNx2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNx2_ASAP7_6t_SL 0 0 ;
  SIZE 1.134 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.176 0.189 ;
        RECT 0.094 0.027 0.176 0.045 ;
        RECT 0.094 0.128 0.117 0.189 ;
        RECT 0.072 0.065 0.115 0.083 ;
        RECT 0.094 0.027 0.115 0.083 ;
        RECT 0.072 0.128 0.117 0.146 ;
        RECT 0.072 0.065 0.09 0.146 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.27 0.027 0.392 0.045 ;
        RECT 0.251 0.171 0.338 0.189 ;
        RECT 0.27 0.027 0.288 0.189 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.951 0.171 1.062 0.189 ;
        RECT 1.044 0.027 1.062 0.189 ;
        RECT 0.951 0.027 1.062 0.045 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.134 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.134 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.881 0.063 0.899 0.126 ;
      RECT 0.862 0.063 0.899 0.081 ;
      RECT 0.81 0.171 0.878 0.189 ;
      RECT 0.81 0.027 0.828 0.189 ;
      RECT 0.769 0.07 0.828 0.088 ;
      RECT 0.809 0.027 0.828 0.088 ;
      RECT 0.809 0.027 0.878 0.045 ;
      RECT 0.688 0.17 0.738 0.188 ;
      RECT 0.72 0.027 0.738 0.188 ;
      RECT 0.634 0.027 0.738 0.045 ;
      RECT 0.666 0.063 0.684 0.123 ;
      RECT 0.654 0.063 0.694 0.081 ;
      RECT 0.601 0.135 0.64 0.153 ;
      RECT 0.612 0.094 0.63 0.153 ;
      RECT 0.522 0.171 0.628 0.189 ;
      RECT 0.522 0.047 0.54 0.189 ;
      RECT 0.494 0.077 0.54 0.095 ;
      RECT 0.522 0.047 0.603 0.065 ;
      RECT 0.369 0.171 0.464 0.189 ;
      RECT 0.446 0.027 0.464 0.189 ;
      RECT 0.423 0.027 0.464 0.045 ;
      RECT 0.396 0.063 0.414 0.126 ;
      RECT 0.377 0.063 0.414 0.081 ;
      RECT 0.306 0.135 0.377 0.153 ;
      RECT 0.306 0.099 0.324 0.153 ;
      RECT 0.306 0.099 0.368 0.117 ;
      RECT 0.201 0.112 0.219 0.158 ;
      RECT 0.201 0.112 0.244 0.13 ;
      RECT 0.225 0.027 0.244 0.13 ;
      RECT 0.207 0.027 0.244 0.045 ;
      RECT 0.143 0.063 0.161 0.117 ;
      RECT 0.143 0.063 0.183 0.081 ;
      RECT 0.016 0.171 0.068 0.189 ;
      RECT 0.016 0.027 0.034 0.189 ;
      RECT 0.016 0.027 0.063 0.045 ;
      RECT 0.774 0.113 0.792 0.172 ;
      RECT 0.558 0.094 0.576 0.144 ;
      RECT 0.486 0.126 0.504 0.172 ;
    LAYER M2 ;
      RECT 0.72 0.063 0.899 0.081 ;
      RECT 0.196 0.135 0.797 0.153 ;
      RECT 0.016 0.063 0.684 0.081 ;
      RECT 0.446 0.099 0.576 0.117 ;
    LAYER V1 ;
      RECT 0.876 0.063 0.894 0.081 ;
      RECT 0.774 0.135 0.792 0.153 ;
      RECT 0.72 0.063 0.738 0.081 ;
      RECT 0.666 0.063 0.684 0.081 ;
      RECT 0.612 0.135 0.63 0.153 ;
      RECT 0.558 0.099 0.576 0.117 ;
      RECT 0.486 0.135 0.504 0.153 ;
      RECT 0.446 0.099 0.464 0.117 ;
      RECT 0.391 0.063 0.409 0.081 ;
      RECT 0.315 0.135 0.333 0.153 ;
      RECT 0.201 0.135 0.219 0.153 ;
      RECT 0.153 0.063 0.171 0.081 ;
      RECT 0.016 0.063 0.034 0.081 ;
  END
END DFFHQNx2_ASAP7_6t_SL

MACRO DFFHQNx3_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNx3_ASAP7_6t_SL 0 0 ;
  SIZE 1.188 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.176 0.189 ;
        RECT 0.094 0.027 0.176 0.045 ;
        RECT 0.094 0.128 0.117 0.189 ;
        RECT 0.072 0.065 0.115 0.083 ;
        RECT 0.094 0.027 0.115 0.083 ;
        RECT 0.072 0.128 0.117 0.146 ;
        RECT 0.072 0.065 0.09 0.146 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.27 0.027 0.392 0.045 ;
        RECT 0.251 0.171 0.338 0.189 ;
        RECT 0.27 0.027 0.288 0.189 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.011 0.171 1.169 0.189 ;
        RECT 1.151 0.027 1.169 0.189 ;
        RECT 1.007 0.027 1.169 0.045 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.188 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.188 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.881 0.063 0.899 0.126 ;
      RECT 0.862 0.063 0.899 0.081 ;
      RECT 0.81 0.171 0.878 0.189 ;
      RECT 0.81 0.027 0.828 0.189 ;
      RECT 0.769 0.07 0.828 0.088 ;
      RECT 0.809 0.027 0.828 0.088 ;
      RECT 0.809 0.027 0.878 0.045 ;
      RECT 0.688 0.17 0.738 0.188 ;
      RECT 0.72 0.027 0.738 0.188 ;
      RECT 0.634 0.027 0.738 0.045 ;
      RECT 0.666 0.063 0.684 0.123 ;
      RECT 0.654 0.063 0.694 0.081 ;
      RECT 0.601 0.135 0.64 0.153 ;
      RECT 0.612 0.094 0.63 0.153 ;
      RECT 0.522 0.171 0.628 0.189 ;
      RECT 0.522 0.047 0.54 0.189 ;
      RECT 0.494 0.077 0.54 0.095 ;
      RECT 0.522 0.047 0.603 0.065 ;
      RECT 0.369 0.171 0.464 0.189 ;
      RECT 0.446 0.027 0.464 0.189 ;
      RECT 0.423 0.027 0.464 0.045 ;
      RECT 0.396 0.063 0.414 0.126 ;
      RECT 0.377 0.063 0.414 0.081 ;
      RECT 0.306 0.135 0.377 0.153 ;
      RECT 0.306 0.099 0.324 0.153 ;
      RECT 0.306 0.099 0.368 0.117 ;
      RECT 0.201 0.112 0.219 0.158 ;
      RECT 0.201 0.112 0.244 0.13 ;
      RECT 0.225 0.027 0.244 0.13 ;
      RECT 0.207 0.027 0.244 0.045 ;
      RECT 0.143 0.063 0.161 0.117 ;
      RECT 0.143 0.063 0.183 0.081 ;
      RECT 0.016 0.171 0.068 0.189 ;
      RECT 0.016 0.027 0.034 0.189 ;
      RECT 0.016 0.027 0.063 0.045 ;
      RECT 0.774 0.113 0.792 0.172 ;
      RECT 0.558 0.094 0.576 0.144 ;
      RECT 0.486 0.126 0.504 0.172 ;
    LAYER M2 ;
      RECT 0.72 0.063 0.899 0.081 ;
      RECT 0.196 0.135 0.797 0.153 ;
      RECT 0.016 0.063 0.684 0.081 ;
      RECT 0.446 0.099 0.576 0.117 ;
    LAYER V1 ;
      RECT 0.876 0.063 0.894 0.081 ;
      RECT 0.774 0.135 0.792 0.153 ;
      RECT 0.72 0.063 0.738 0.081 ;
      RECT 0.666 0.063 0.684 0.081 ;
      RECT 0.612 0.135 0.63 0.153 ;
      RECT 0.558 0.099 0.576 0.117 ;
      RECT 0.486 0.135 0.504 0.153 ;
      RECT 0.446 0.099 0.464 0.117 ;
      RECT 0.391 0.063 0.409 0.081 ;
      RECT 0.315 0.135 0.333 0.153 ;
      RECT 0.201 0.135 0.219 0.153 ;
      RECT 0.153 0.063 0.171 0.081 ;
      RECT 0.016 0.063 0.034 0.081 ;
  END
END DFFHQNx3_ASAP7_6t_SL

MACRO DFFHQx4_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQx4_ASAP7_6t_SL 0 0 ;
  SIZE 1.35 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.176 0.189 ;
        RECT 0.094 0.027 0.176 0.045 ;
        RECT 0.094 0.128 0.117 0.189 ;
        RECT 0.072 0.065 0.115 0.083 ;
        RECT 0.094 0.027 0.115 0.083 ;
        RECT 0.072 0.128 0.117 0.146 ;
        RECT 0.072 0.065 0.09 0.146 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.27 0.027 0.392 0.045 ;
        RECT 0.251 0.171 0.338 0.189 ;
        RECT 0.27 0.027 0.288 0.189 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.125 0.171 1.333 0.189 ;
        RECT 1.313 0.027 1.333 0.189 ;
        RECT 1.125 0.027 1.333 0.045 ;
        RECT 1.125 0.147 1.143 0.189 ;
        RECT 1.125 0.027 1.143 0.069 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.35 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.35 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.012 0.171 1.098 0.189 ;
      RECT 1.08 0.027 1.098 0.189 ;
      RECT 1.08 0.1 1.175 0.118 ;
      RECT 1.012 0.027 1.098 0.045 ;
      RECT 0.881 0.063 0.899 0.126 ;
      RECT 0.862 0.063 0.899 0.081 ;
      RECT 0.81 0.171 0.878 0.189 ;
      RECT 0.81 0.027 0.828 0.189 ;
      RECT 0.769 0.07 0.828 0.088 ;
      RECT 0.809 0.027 0.828 0.088 ;
      RECT 0.809 0.027 0.878 0.045 ;
      RECT 0.688 0.17 0.738 0.188 ;
      RECT 0.72 0.027 0.738 0.188 ;
      RECT 0.634 0.027 0.738 0.045 ;
      RECT 0.666 0.063 0.684 0.123 ;
      RECT 0.654 0.063 0.694 0.081 ;
      RECT 0.601 0.135 0.64 0.153 ;
      RECT 0.612 0.094 0.63 0.153 ;
      RECT 0.522 0.171 0.628 0.189 ;
      RECT 0.522 0.047 0.54 0.189 ;
      RECT 0.494 0.077 0.54 0.095 ;
      RECT 0.522 0.047 0.603 0.065 ;
      RECT 0.369 0.171 0.464 0.189 ;
      RECT 0.446 0.027 0.464 0.189 ;
      RECT 0.423 0.027 0.464 0.045 ;
      RECT 0.396 0.063 0.414 0.126 ;
      RECT 0.377 0.063 0.414 0.081 ;
      RECT 0.306 0.135 0.377 0.153 ;
      RECT 0.306 0.099 0.324 0.153 ;
      RECT 0.306 0.099 0.368 0.117 ;
      RECT 0.201 0.112 0.219 0.158 ;
      RECT 0.201 0.112 0.244 0.13 ;
      RECT 0.225 0.027 0.244 0.13 ;
      RECT 0.207 0.027 0.244 0.045 ;
      RECT 0.143 0.063 0.161 0.117 ;
      RECT 0.143 0.063 0.183 0.081 ;
      RECT 0.016 0.171 0.068 0.189 ;
      RECT 0.016 0.027 0.034 0.189 ;
      RECT 0.016 0.027 0.063 0.045 ;
      RECT 0.774 0.113 0.792 0.172 ;
      RECT 0.558 0.094 0.576 0.144 ;
      RECT 0.486 0.126 0.504 0.172 ;
    LAYER M2 ;
      RECT 0.72 0.063 0.899 0.081 ;
      RECT 0.196 0.135 0.797 0.153 ;
      RECT 0.016 0.063 0.684 0.081 ;
      RECT 0.446 0.099 0.576 0.117 ;
    LAYER V1 ;
      RECT 0.876 0.063 0.894 0.081 ;
      RECT 0.774 0.135 0.792 0.153 ;
      RECT 0.72 0.063 0.738 0.081 ;
      RECT 0.666 0.063 0.684 0.081 ;
      RECT 0.612 0.135 0.63 0.153 ;
      RECT 0.558 0.099 0.576 0.117 ;
      RECT 0.486 0.135 0.504 0.153 ;
      RECT 0.446 0.099 0.464 0.117 ;
      RECT 0.391 0.063 0.409 0.081 ;
      RECT 0.315 0.135 0.333 0.153 ;
      RECT 0.201 0.135 0.219 0.153 ;
      RECT 0.153 0.063 0.171 0.081 ;
      RECT 0.016 0.063 0.034 0.081 ;
  END
END DFFHQx4_ASAP7_6t_SL

MACRO DFFLQNx1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFLQNx1_ASAP7_6t_SL 0 0 ;
  SIZE 1.08 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.176 0.189 ;
        RECT 0.094 0.027 0.176 0.045 ;
        RECT 0.072 0.07 0.117 0.088 ;
        RECT 0.094 0.027 0.117 0.088 ;
        RECT 0.094 0.133 0.115 0.189 ;
        RECT 0.072 0.133 0.115 0.151 ;
        RECT 0.072 0.07 0.09 0.151 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.27 0.171 0.392 0.189 ;
        RECT 0.251 0.027 0.338 0.045 ;
        RECT 0.27 0.027 0.288 0.189 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.953 0.171 1.062 0.189 ;
        RECT 1.044 0.027 1.062 0.189 ;
        RECT 0.953 0.027 1.062 0.045 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.08 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.08 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.862 0.135 0.899 0.153 ;
      RECT 0.881 0.09 0.899 0.153 ;
      RECT 0.809 0.171 0.878 0.189 ;
      RECT 0.809 0.128 0.828 0.189 ;
      RECT 0.81 0.027 0.828 0.189 ;
      RECT 0.769 0.128 0.828 0.146 ;
      RECT 0.81 0.027 0.878 0.045 ;
      RECT 0.634 0.171 0.738 0.189 ;
      RECT 0.72 0.028 0.738 0.189 ;
      RECT 0.688 0.028 0.738 0.046 ;
      RECT 0.654 0.135 0.694 0.153 ;
      RECT 0.666 0.093 0.684 0.153 ;
      RECT 0.612 0.063 0.63 0.122 ;
      RECT 0.601 0.063 0.64 0.081 ;
      RECT 0.522 0.151 0.603 0.169 ;
      RECT 0.522 0.027 0.54 0.169 ;
      RECT 0.494 0.121 0.54 0.139 ;
      RECT 0.522 0.027 0.628 0.045 ;
      RECT 0.423 0.171 0.464 0.189 ;
      RECT 0.446 0.027 0.464 0.189 ;
      RECT 0.369 0.027 0.464 0.045 ;
      RECT 0.377 0.135 0.414 0.153 ;
      RECT 0.396 0.09 0.414 0.153 ;
      RECT 0.306 0.099 0.368 0.117 ;
      RECT 0.306 0.063 0.324 0.117 ;
      RECT 0.306 0.063 0.377 0.081 ;
      RECT 0.207 0.171 0.244 0.189 ;
      RECT 0.225 0.086 0.244 0.189 ;
      RECT 0.201 0.086 0.244 0.104 ;
      RECT 0.201 0.058 0.219 0.104 ;
      RECT 0.143 0.135 0.183 0.153 ;
      RECT 0.143 0.099 0.161 0.153 ;
      RECT 0.016 0.171 0.063 0.189 ;
      RECT 0.016 0.027 0.034 0.189 ;
      RECT 0.016 0.027 0.068 0.045 ;
      RECT 0.774 0.044 0.792 0.103 ;
      RECT 0.558 0.072 0.576 0.122 ;
      RECT 0.486 0.044 0.504 0.09 ;
    LAYER M2 ;
      RECT 0.72 0.135 0.899 0.153 ;
      RECT 0.196 0.063 0.797 0.081 ;
      RECT 0.016 0.135 0.684 0.153 ;
      RECT 0.446 0.099 0.576 0.117 ;
    LAYER V1 ;
      RECT 0.876 0.135 0.894 0.153 ;
      RECT 0.774 0.063 0.792 0.081 ;
      RECT 0.72 0.135 0.738 0.153 ;
      RECT 0.666 0.135 0.684 0.153 ;
      RECT 0.612 0.063 0.63 0.081 ;
      RECT 0.558 0.099 0.576 0.117 ;
      RECT 0.486 0.063 0.504 0.081 ;
      RECT 0.446 0.099 0.464 0.117 ;
      RECT 0.391 0.135 0.409 0.153 ;
      RECT 0.315 0.063 0.333 0.081 ;
      RECT 0.201 0.063 0.219 0.081 ;
      RECT 0.153 0.135 0.171 0.153 ;
      RECT 0.016 0.135 0.034 0.153 ;
  END
END DFFLQNx1_ASAP7_6t_SL

MACRO DFFLQNx2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFLQNx2_ASAP7_6t_SL 0 0 ;
  SIZE 1.134 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.176 0.189 ;
        RECT 0.094 0.027 0.176 0.045 ;
        RECT 0.072 0.07 0.117 0.088 ;
        RECT 0.094 0.027 0.117 0.088 ;
        RECT 0.094 0.133 0.115 0.189 ;
        RECT 0.072 0.133 0.115 0.151 ;
        RECT 0.072 0.07 0.09 0.151 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.27 0.171 0.392 0.189 ;
        RECT 0.251 0.027 0.338 0.045 ;
        RECT 0.27 0.027 0.288 0.189 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.953 0.171 1.062 0.189 ;
        RECT 1.044 0.027 1.062 0.189 ;
        RECT 0.953 0.027 1.062 0.045 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.134 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.134 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.862 0.135 0.899 0.153 ;
      RECT 0.881 0.09 0.899 0.153 ;
      RECT 0.809 0.171 0.878 0.189 ;
      RECT 0.809 0.128 0.828 0.189 ;
      RECT 0.81 0.027 0.828 0.189 ;
      RECT 0.769 0.128 0.828 0.146 ;
      RECT 0.81 0.027 0.878 0.045 ;
      RECT 0.634 0.171 0.738 0.189 ;
      RECT 0.72 0.028 0.738 0.189 ;
      RECT 0.688 0.028 0.738 0.046 ;
      RECT 0.654 0.135 0.694 0.153 ;
      RECT 0.666 0.093 0.684 0.153 ;
      RECT 0.612 0.063 0.63 0.122 ;
      RECT 0.601 0.063 0.64 0.081 ;
      RECT 0.522 0.151 0.603 0.169 ;
      RECT 0.522 0.027 0.54 0.169 ;
      RECT 0.494 0.121 0.54 0.139 ;
      RECT 0.522 0.027 0.628 0.045 ;
      RECT 0.423 0.171 0.464 0.189 ;
      RECT 0.446 0.027 0.464 0.189 ;
      RECT 0.369 0.027 0.464 0.045 ;
      RECT 0.377 0.135 0.414 0.153 ;
      RECT 0.396 0.09 0.414 0.153 ;
      RECT 0.306 0.099 0.368 0.117 ;
      RECT 0.306 0.063 0.324 0.117 ;
      RECT 0.306 0.063 0.377 0.081 ;
      RECT 0.207 0.171 0.244 0.189 ;
      RECT 0.225 0.086 0.244 0.189 ;
      RECT 0.201 0.086 0.244 0.104 ;
      RECT 0.201 0.058 0.219 0.104 ;
      RECT 0.143 0.135 0.183 0.153 ;
      RECT 0.143 0.099 0.161 0.153 ;
      RECT 0.016 0.171 0.063 0.189 ;
      RECT 0.016 0.027 0.034 0.189 ;
      RECT 0.016 0.027 0.068 0.045 ;
      RECT 0.774 0.044 0.792 0.103 ;
      RECT 0.558 0.072 0.576 0.122 ;
      RECT 0.486 0.044 0.504 0.09 ;
    LAYER M2 ;
      RECT 0.72 0.135 0.899 0.153 ;
      RECT 0.196 0.063 0.797 0.081 ;
      RECT 0.016 0.135 0.684 0.153 ;
      RECT 0.446 0.099 0.576 0.117 ;
    LAYER V1 ;
      RECT 0.876 0.135 0.894 0.153 ;
      RECT 0.774 0.063 0.792 0.081 ;
      RECT 0.72 0.135 0.738 0.153 ;
      RECT 0.666 0.135 0.684 0.153 ;
      RECT 0.612 0.063 0.63 0.081 ;
      RECT 0.558 0.099 0.576 0.117 ;
      RECT 0.486 0.063 0.504 0.081 ;
      RECT 0.446 0.099 0.464 0.117 ;
      RECT 0.391 0.135 0.409 0.153 ;
      RECT 0.315 0.063 0.333 0.081 ;
      RECT 0.201 0.063 0.219 0.081 ;
      RECT 0.153 0.135 0.171 0.153 ;
      RECT 0.016 0.135 0.034 0.153 ;
  END
END DFFLQNx2_ASAP7_6t_SL

MACRO DFFLQNx3_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFLQNx3_ASAP7_6t_SL 0 0 ;
  SIZE 1.188 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.176 0.189 ;
        RECT 0.094 0.027 0.176 0.045 ;
        RECT 0.072 0.07 0.117 0.088 ;
        RECT 0.094 0.027 0.117 0.088 ;
        RECT 0.094 0.133 0.115 0.189 ;
        RECT 0.072 0.133 0.115 0.151 ;
        RECT 0.072 0.07 0.09 0.151 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.27 0.171 0.392 0.189 ;
        RECT 0.251 0.027 0.338 0.045 ;
        RECT 0.27 0.027 0.288 0.189 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.007 0.171 1.169 0.189 ;
        RECT 1.151 0.027 1.169 0.189 ;
        RECT 1.011 0.027 1.169 0.045 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.188 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.188 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.862 0.135 0.899 0.153 ;
      RECT 0.881 0.09 0.899 0.153 ;
      RECT 0.809 0.171 0.878 0.189 ;
      RECT 0.809 0.128 0.828 0.189 ;
      RECT 0.81 0.027 0.828 0.189 ;
      RECT 0.769 0.128 0.828 0.146 ;
      RECT 0.81 0.027 0.878 0.045 ;
      RECT 0.634 0.171 0.738 0.189 ;
      RECT 0.72 0.028 0.738 0.189 ;
      RECT 0.688 0.028 0.738 0.046 ;
      RECT 0.654 0.135 0.694 0.153 ;
      RECT 0.666 0.093 0.684 0.153 ;
      RECT 0.612 0.063 0.63 0.122 ;
      RECT 0.601 0.063 0.64 0.081 ;
      RECT 0.522 0.151 0.603 0.169 ;
      RECT 0.522 0.027 0.54 0.169 ;
      RECT 0.494 0.121 0.54 0.139 ;
      RECT 0.522 0.027 0.628 0.045 ;
      RECT 0.423 0.171 0.464 0.189 ;
      RECT 0.446 0.027 0.464 0.189 ;
      RECT 0.369 0.027 0.464 0.045 ;
      RECT 0.377 0.135 0.414 0.153 ;
      RECT 0.396 0.09 0.414 0.153 ;
      RECT 0.306 0.099 0.368 0.117 ;
      RECT 0.306 0.063 0.324 0.117 ;
      RECT 0.306 0.063 0.377 0.081 ;
      RECT 0.207 0.171 0.244 0.189 ;
      RECT 0.225 0.086 0.244 0.189 ;
      RECT 0.201 0.086 0.244 0.104 ;
      RECT 0.201 0.058 0.219 0.104 ;
      RECT 0.143 0.135 0.183 0.153 ;
      RECT 0.143 0.099 0.161 0.153 ;
      RECT 0.016 0.171 0.063 0.189 ;
      RECT 0.016 0.027 0.034 0.189 ;
      RECT 0.016 0.027 0.068 0.045 ;
      RECT 0.774 0.044 0.792 0.103 ;
      RECT 0.558 0.072 0.576 0.122 ;
      RECT 0.486 0.044 0.504 0.09 ;
    LAYER M2 ;
      RECT 0.72 0.135 0.899 0.153 ;
      RECT 0.196 0.063 0.797 0.081 ;
      RECT 0.016 0.135 0.684 0.153 ;
      RECT 0.446 0.099 0.576 0.117 ;
    LAYER V1 ;
      RECT 0.876 0.135 0.894 0.153 ;
      RECT 0.774 0.063 0.792 0.081 ;
      RECT 0.72 0.135 0.738 0.153 ;
      RECT 0.666 0.135 0.684 0.153 ;
      RECT 0.612 0.063 0.63 0.081 ;
      RECT 0.558 0.099 0.576 0.117 ;
      RECT 0.486 0.063 0.504 0.081 ;
      RECT 0.446 0.099 0.464 0.117 ;
      RECT 0.391 0.135 0.409 0.153 ;
      RECT 0.315 0.063 0.333 0.081 ;
      RECT 0.201 0.063 0.219 0.081 ;
      RECT 0.153 0.135 0.171 0.153 ;
      RECT 0.016 0.135 0.034 0.153 ;
  END
END DFFLQNx3_ASAP7_6t_SL

MACRO DFFLQx4_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFLQx4_ASAP7_6t_SL 0 0 ;
  SIZE 1.35 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.176 0.189 ;
        RECT 0.094 0.027 0.176 0.045 ;
        RECT 0.072 0.07 0.117 0.088 ;
        RECT 0.094 0.027 0.117 0.088 ;
        RECT 0.094 0.133 0.115 0.189 ;
        RECT 0.072 0.133 0.115 0.151 ;
        RECT 0.072 0.07 0.09 0.151 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.27 0.171 0.392 0.189 ;
        RECT 0.251 0.027 0.338 0.045 ;
        RECT 0.27 0.027 0.288 0.189 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.125 0.171 1.333 0.189 ;
        RECT 1.313 0.027 1.333 0.189 ;
        RECT 1.125 0.027 1.333 0.045 ;
        RECT 1.125 0.147 1.143 0.189 ;
        RECT 1.125 0.027 1.143 0.069 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.35 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.35 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.012 0.171 1.098 0.189 ;
      RECT 1.08 0.027 1.098 0.189 ;
      RECT 1.08 0.098 1.175 0.116 ;
      RECT 1.012 0.027 1.098 0.045 ;
      RECT 0.862 0.135 0.899 0.153 ;
      RECT 0.881 0.09 0.899 0.153 ;
      RECT 0.809 0.171 0.878 0.189 ;
      RECT 0.809 0.128 0.828 0.189 ;
      RECT 0.81 0.027 0.828 0.189 ;
      RECT 0.769 0.128 0.828 0.146 ;
      RECT 0.81 0.027 0.878 0.045 ;
      RECT 0.634 0.171 0.738 0.189 ;
      RECT 0.72 0.028 0.738 0.189 ;
      RECT 0.688 0.028 0.738 0.046 ;
      RECT 0.654 0.135 0.694 0.153 ;
      RECT 0.666 0.093 0.684 0.153 ;
      RECT 0.612 0.063 0.63 0.122 ;
      RECT 0.601 0.063 0.64 0.081 ;
      RECT 0.522 0.151 0.603 0.169 ;
      RECT 0.522 0.027 0.54 0.169 ;
      RECT 0.494 0.121 0.54 0.139 ;
      RECT 0.522 0.027 0.628 0.045 ;
      RECT 0.423 0.171 0.464 0.189 ;
      RECT 0.446 0.027 0.464 0.189 ;
      RECT 0.369 0.027 0.464 0.045 ;
      RECT 0.377 0.135 0.414 0.153 ;
      RECT 0.396 0.09 0.414 0.153 ;
      RECT 0.306 0.099 0.368 0.117 ;
      RECT 0.306 0.063 0.324 0.117 ;
      RECT 0.306 0.063 0.377 0.081 ;
      RECT 0.207 0.171 0.244 0.189 ;
      RECT 0.225 0.086 0.244 0.189 ;
      RECT 0.201 0.086 0.244 0.104 ;
      RECT 0.201 0.058 0.219 0.104 ;
      RECT 0.143 0.135 0.183 0.153 ;
      RECT 0.143 0.099 0.161 0.153 ;
      RECT 0.016 0.171 0.063 0.189 ;
      RECT 0.016 0.027 0.034 0.189 ;
      RECT 0.016 0.027 0.068 0.045 ;
      RECT 0.774 0.044 0.792 0.103 ;
      RECT 0.558 0.072 0.576 0.122 ;
      RECT 0.486 0.044 0.504 0.09 ;
    LAYER M2 ;
      RECT 0.72 0.135 0.899 0.153 ;
      RECT 0.196 0.063 0.797 0.081 ;
      RECT 0.016 0.135 0.684 0.153 ;
      RECT 0.446 0.099 0.576 0.117 ;
    LAYER V1 ;
      RECT 0.876 0.135 0.894 0.153 ;
      RECT 0.774 0.063 0.792 0.081 ;
      RECT 0.72 0.135 0.738 0.153 ;
      RECT 0.666 0.135 0.684 0.153 ;
      RECT 0.612 0.063 0.63 0.081 ;
      RECT 0.558 0.099 0.576 0.117 ;
      RECT 0.486 0.063 0.504 0.081 ;
      RECT 0.446 0.099 0.464 0.117 ;
      RECT 0.391 0.135 0.409 0.153 ;
      RECT 0.315 0.063 0.333 0.081 ;
      RECT 0.201 0.063 0.219 0.081 ;
      RECT 0.153 0.135 0.171 0.153 ;
      RECT 0.016 0.135 0.034 0.153 ;
  END
END DFFLQx4_ASAP7_6t_SL

MACRO DHLx1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHLx1_ASAP7_6t_SL 0 0 ;
  SIZE 0.81 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.176 0.189 ;
        RECT 0.094 0.027 0.176 0.045 ;
        RECT 0.072 0.065 0.117 0.083 ;
        RECT 0.094 0.027 0.117 0.083 ;
        RECT 0.094 0.128 0.112 0.189 ;
        RECT 0.072 0.128 0.112 0.146 ;
        RECT 0.072 0.065 0.09 0.146 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.27 0.171 0.338 0.189 ;
        RECT 0.27 0.027 0.338 0.045 ;
        RECT 0.27 0.099 0.306 0.117 ;
        RECT 0.27 0.027 0.288 0.189 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.686 0.171 0.792 0.189 ;
        RECT 0.774 0.027 0.792 0.189 ;
        RECT 0.686 0.027 0.792 0.045 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.81 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.81 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.58 0.171 0.657 0.189 ;
      RECT 0.639 0.027 0.657 0.189 ;
      RECT 0.504 0.07 0.552 0.088 ;
      RECT 0.534 0.027 0.552 0.088 ;
      RECT 0.534 0.027 0.657 0.045 ;
      RECT 0.603 0.063 0.621 0.126 ;
      RECT 0.577 0.063 0.621 0.081 ;
      RECT 0.369 0.171 0.468 0.189 ;
      RECT 0.45 0.027 0.468 0.189 ;
      RECT 0.413 0.027 0.468 0.045 ;
      RECT 0.396 0.063 0.414 0.126 ;
      RECT 0.382 0.063 0.424 0.081 ;
      RECT 0.338 0.135 0.375 0.153 ;
      RECT 0.342 0.085 0.36 0.153 ;
      RECT 0.207 0.171 0.245 0.189 ;
      RECT 0.227 0.027 0.245 0.189 ;
      RECT 0.207 0.027 0.245 0.045 ;
      RECT 0.143 0.135 0.198 0.153 ;
      RECT 0.18 0.099 0.198 0.153 ;
      RECT 0.138 0.099 0.198 0.117 ;
      RECT 0.016 0.171 0.068 0.189 ;
      RECT 0.016 0.027 0.034 0.189 ;
      RECT 0.016 0.027 0.068 0.045 ;
      RECT 0.504 0.113 0.522 0.172 ;
    LAYER M2 ;
      RECT 0.45 0.063 0.61 0.081 ;
      RECT 0.016 0.135 0.527 0.153 ;
      RECT 0.222 0.063 0.414 0.081 ;
    LAYER V1 ;
      RECT 0.585 0.063 0.603 0.081 ;
      RECT 0.504 0.135 0.522 0.153 ;
      RECT 0.45 0.063 0.468 0.081 ;
      RECT 0.396 0.063 0.414 0.081 ;
      RECT 0.342 0.135 0.36 0.153 ;
      RECT 0.227 0.063 0.245 0.081 ;
      RECT 0.153 0.135 0.171 0.153 ;
      RECT 0.016 0.135 0.034 0.153 ;
  END
END DHLx1_ASAP7_6t_SL

MACRO DHLx2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHLx2_ASAP7_6t_SL 0 0 ;
  SIZE 0.864 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.176 0.189 ;
        RECT 0.094 0.027 0.176 0.045 ;
        RECT 0.072 0.065 0.117 0.083 ;
        RECT 0.094 0.027 0.117 0.083 ;
        RECT 0.094 0.128 0.112 0.189 ;
        RECT 0.072 0.128 0.112 0.146 ;
        RECT 0.072 0.065 0.09 0.146 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.27 0.171 0.338 0.189 ;
        RECT 0.27 0.027 0.338 0.045 ;
        RECT 0.27 0.099 0.306 0.117 ;
        RECT 0.27 0.027 0.288 0.189 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.688 0.171 0.792 0.189 ;
        RECT 0.774 0.027 0.792 0.189 ;
        RECT 0.688 0.027 0.792 0.045 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.864 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.864 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.58 0.171 0.657 0.189 ;
      RECT 0.639 0.027 0.657 0.189 ;
      RECT 0.504 0.07 0.552 0.088 ;
      RECT 0.534 0.027 0.552 0.088 ;
      RECT 0.534 0.027 0.657 0.045 ;
      RECT 0.603 0.063 0.621 0.126 ;
      RECT 0.577 0.063 0.621 0.081 ;
      RECT 0.369 0.171 0.468 0.189 ;
      RECT 0.45 0.027 0.468 0.189 ;
      RECT 0.413 0.027 0.468 0.045 ;
      RECT 0.396 0.063 0.414 0.126 ;
      RECT 0.382 0.063 0.424 0.081 ;
      RECT 0.338 0.135 0.375 0.153 ;
      RECT 0.342 0.085 0.36 0.153 ;
      RECT 0.207 0.171 0.245 0.189 ;
      RECT 0.227 0.027 0.245 0.189 ;
      RECT 0.207 0.027 0.245 0.045 ;
      RECT 0.143 0.135 0.198 0.153 ;
      RECT 0.18 0.099 0.198 0.153 ;
      RECT 0.138 0.099 0.198 0.117 ;
      RECT 0.016 0.171 0.068 0.189 ;
      RECT 0.016 0.027 0.034 0.189 ;
      RECT 0.016 0.027 0.068 0.045 ;
      RECT 0.504 0.113 0.522 0.172 ;
    LAYER M2 ;
      RECT 0.45 0.063 0.61 0.081 ;
      RECT 0.016 0.135 0.527 0.153 ;
      RECT 0.222 0.063 0.414 0.081 ;
    LAYER V1 ;
      RECT 0.585 0.063 0.603 0.081 ;
      RECT 0.504 0.135 0.522 0.153 ;
      RECT 0.45 0.063 0.468 0.081 ;
      RECT 0.396 0.063 0.414 0.081 ;
      RECT 0.342 0.135 0.36 0.153 ;
      RECT 0.227 0.063 0.245 0.081 ;
      RECT 0.153 0.135 0.171 0.153 ;
      RECT 0.016 0.135 0.034 0.153 ;
  END
END DHLx2_ASAP7_6t_SL

MACRO DHLx3_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHLx3_ASAP7_6t_SL 0 0 ;
  SIZE 0.918 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.176 0.189 ;
        RECT 0.094 0.027 0.176 0.045 ;
        RECT 0.072 0.065 0.117 0.083 ;
        RECT 0.094 0.027 0.117 0.083 ;
        RECT 0.094 0.128 0.112 0.189 ;
        RECT 0.072 0.128 0.112 0.146 ;
        RECT 0.072 0.065 0.09 0.146 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.27 0.171 0.338 0.189 ;
        RECT 0.27 0.027 0.338 0.045 ;
        RECT 0.27 0.099 0.306 0.117 ;
        RECT 0.27 0.027 0.288 0.189 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.724 0.171 0.881 0.189 ;
        RECT 0.727 0.027 0.881 0.045 ;
        RECT 0.774 0.027 0.792 0.189 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.918 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.918 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.58 0.171 0.657 0.189 ;
      RECT 0.639 0.027 0.657 0.189 ;
      RECT 0.504 0.07 0.552 0.088 ;
      RECT 0.534 0.027 0.552 0.088 ;
      RECT 0.534 0.027 0.657 0.045 ;
      RECT 0.603 0.063 0.621 0.126 ;
      RECT 0.577 0.063 0.621 0.081 ;
      RECT 0.369 0.171 0.468 0.189 ;
      RECT 0.45 0.027 0.468 0.189 ;
      RECT 0.413 0.027 0.468 0.045 ;
      RECT 0.396 0.063 0.414 0.126 ;
      RECT 0.382 0.063 0.424 0.081 ;
      RECT 0.338 0.135 0.375 0.153 ;
      RECT 0.342 0.085 0.36 0.153 ;
      RECT 0.207 0.171 0.245 0.189 ;
      RECT 0.227 0.027 0.245 0.189 ;
      RECT 0.207 0.027 0.245 0.045 ;
      RECT 0.143 0.135 0.198 0.153 ;
      RECT 0.18 0.099 0.198 0.153 ;
      RECT 0.138 0.099 0.198 0.117 ;
      RECT 0.016 0.171 0.068 0.189 ;
      RECT 0.016 0.027 0.034 0.189 ;
      RECT 0.016 0.027 0.068 0.045 ;
      RECT 0.504 0.113 0.522 0.172 ;
    LAYER M2 ;
      RECT 0.45 0.063 0.61 0.081 ;
      RECT 0.016 0.135 0.527 0.153 ;
      RECT 0.222 0.063 0.414 0.081 ;
    LAYER V1 ;
      RECT 0.585 0.063 0.603 0.081 ;
      RECT 0.504 0.135 0.522 0.153 ;
      RECT 0.45 0.063 0.468 0.081 ;
      RECT 0.396 0.063 0.414 0.081 ;
      RECT 0.342 0.135 0.36 0.153 ;
      RECT 0.227 0.063 0.245 0.081 ;
      RECT 0.153 0.135 0.171 0.153 ;
      RECT 0.016 0.135 0.034 0.153 ;
  END
END DHLx3_ASAP7_6t_SL

MACRO DLLx1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLLx1_ASAP7_6t_SL 0 0 ;
  SIZE 0.81 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.176 0.189 ;
        RECT 0.094 0.027 0.176 0.045 ;
        RECT 0.094 0.133 0.117 0.189 ;
        RECT 0.072 0.07 0.112 0.088 ;
        RECT 0.094 0.027 0.112 0.088 ;
        RECT 0.072 0.133 0.117 0.151 ;
        RECT 0.072 0.07 0.09 0.151 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.27 0.171 0.338 0.189 ;
        RECT 0.27 0.027 0.338 0.045 ;
        RECT 0.27 0.099 0.306 0.117 ;
        RECT 0.27 0.027 0.288 0.189 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.686 0.171 0.792 0.189 ;
        RECT 0.774 0.027 0.792 0.189 ;
        RECT 0.686 0.027 0.792 0.045 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.81 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.81 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.534 0.171 0.657 0.189 ;
      RECT 0.639 0.027 0.657 0.189 ;
      RECT 0.534 0.128 0.552 0.189 ;
      RECT 0.504 0.128 0.552 0.146 ;
      RECT 0.58 0.027 0.657 0.045 ;
      RECT 0.577 0.135 0.621 0.153 ;
      RECT 0.603 0.09 0.621 0.153 ;
      RECT 0.413 0.171 0.468 0.189 ;
      RECT 0.45 0.027 0.468 0.189 ;
      RECT 0.369 0.027 0.468 0.045 ;
      RECT 0.382 0.135 0.424 0.153 ;
      RECT 0.396 0.09 0.414 0.153 ;
      RECT 0.342 0.063 0.36 0.131 ;
      RECT 0.338 0.063 0.375 0.081 ;
      RECT 0.207 0.171 0.245 0.189 ;
      RECT 0.227 0.027 0.245 0.189 ;
      RECT 0.207 0.027 0.245 0.045 ;
      RECT 0.138 0.099 0.198 0.117 ;
      RECT 0.18 0.063 0.198 0.117 ;
      RECT 0.143 0.063 0.198 0.081 ;
      RECT 0.016 0.171 0.068 0.189 ;
      RECT 0.016 0.027 0.034 0.189 ;
      RECT 0.016 0.027 0.068 0.045 ;
      RECT 0.504 0.044 0.522 0.103 ;
    LAYER M2 ;
      RECT 0.45 0.135 0.61 0.153 ;
      RECT 0.016 0.063 0.527 0.081 ;
      RECT 0.222 0.135 0.414 0.153 ;
    LAYER V1 ;
      RECT 0.585 0.135 0.603 0.153 ;
      RECT 0.504 0.063 0.522 0.081 ;
      RECT 0.45 0.135 0.468 0.153 ;
      RECT 0.396 0.135 0.414 0.153 ;
      RECT 0.342 0.063 0.36 0.081 ;
      RECT 0.227 0.135 0.245 0.153 ;
      RECT 0.153 0.063 0.171 0.081 ;
      RECT 0.016 0.063 0.034 0.081 ;
  END
END DLLx1_ASAP7_6t_SL

MACRO DLLx2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLLx2_ASAP7_6t_SL 0 0 ;
  SIZE 0.864 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.176 0.189 ;
        RECT 0.094 0.027 0.176 0.045 ;
        RECT 0.094 0.133 0.117 0.189 ;
        RECT 0.072 0.07 0.112 0.088 ;
        RECT 0.094 0.027 0.112 0.088 ;
        RECT 0.072 0.133 0.117 0.151 ;
        RECT 0.072 0.07 0.09 0.151 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.27 0.171 0.338 0.189 ;
        RECT 0.27 0.027 0.338 0.045 ;
        RECT 0.27 0.099 0.306 0.117 ;
        RECT 0.27 0.027 0.288 0.189 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.686 0.171 0.792 0.189 ;
        RECT 0.774 0.027 0.792 0.189 ;
        RECT 0.686 0.027 0.792 0.045 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.864 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.864 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.534 0.171 0.657 0.189 ;
      RECT 0.639 0.027 0.657 0.189 ;
      RECT 0.534 0.128 0.552 0.189 ;
      RECT 0.504 0.128 0.552 0.146 ;
      RECT 0.58 0.027 0.657 0.045 ;
      RECT 0.577 0.135 0.621 0.153 ;
      RECT 0.603 0.09 0.621 0.153 ;
      RECT 0.413 0.171 0.468 0.189 ;
      RECT 0.45 0.027 0.468 0.189 ;
      RECT 0.369 0.027 0.468 0.045 ;
      RECT 0.382 0.135 0.424 0.153 ;
      RECT 0.396 0.09 0.414 0.153 ;
      RECT 0.342 0.063 0.36 0.131 ;
      RECT 0.338 0.063 0.375 0.081 ;
      RECT 0.207 0.171 0.245 0.189 ;
      RECT 0.227 0.027 0.245 0.189 ;
      RECT 0.207 0.027 0.245 0.045 ;
      RECT 0.138 0.099 0.198 0.117 ;
      RECT 0.18 0.063 0.198 0.117 ;
      RECT 0.143 0.063 0.198 0.081 ;
      RECT 0.016 0.171 0.068 0.189 ;
      RECT 0.016 0.027 0.034 0.189 ;
      RECT 0.016 0.027 0.068 0.045 ;
      RECT 0.504 0.044 0.522 0.103 ;
    LAYER M2 ;
      RECT 0.45 0.135 0.61 0.153 ;
      RECT 0.016 0.063 0.527 0.081 ;
      RECT 0.222 0.135 0.414 0.153 ;
    LAYER V1 ;
      RECT 0.585 0.135 0.603 0.153 ;
      RECT 0.504 0.063 0.522 0.081 ;
      RECT 0.45 0.135 0.468 0.153 ;
      RECT 0.396 0.135 0.414 0.153 ;
      RECT 0.342 0.063 0.36 0.081 ;
      RECT 0.227 0.135 0.245 0.153 ;
      RECT 0.153 0.063 0.171 0.081 ;
      RECT 0.016 0.063 0.034 0.081 ;
  END
END DLLx2_ASAP7_6t_SL

MACRO DLLx3_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLLx3_ASAP7_6t_SL 0 0 ;
  SIZE 0.918 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.176 0.189 ;
        RECT 0.094 0.027 0.176 0.045 ;
        RECT 0.094 0.133 0.117 0.189 ;
        RECT 0.072 0.07 0.112 0.088 ;
        RECT 0.094 0.027 0.112 0.088 ;
        RECT 0.072 0.133 0.117 0.151 ;
        RECT 0.072 0.07 0.09 0.151 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.27 0.171 0.338 0.189 ;
        RECT 0.27 0.027 0.338 0.045 ;
        RECT 0.27 0.099 0.306 0.117 ;
        RECT 0.27 0.027 0.288 0.189 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.727 0.171 0.881 0.189 ;
        RECT 0.723 0.027 0.881 0.045 ;
        RECT 0.774 0.027 0.792 0.189 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.918 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.918 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.534 0.171 0.657 0.189 ;
      RECT 0.639 0.027 0.657 0.189 ;
      RECT 0.534 0.128 0.552 0.189 ;
      RECT 0.504 0.128 0.552 0.146 ;
      RECT 0.58 0.027 0.657 0.045 ;
      RECT 0.577 0.135 0.621 0.153 ;
      RECT 0.603 0.09 0.621 0.153 ;
      RECT 0.413 0.171 0.468 0.189 ;
      RECT 0.45 0.027 0.468 0.189 ;
      RECT 0.369 0.027 0.468 0.045 ;
      RECT 0.382 0.135 0.424 0.153 ;
      RECT 0.396 0.09 0.414 0.153 ;
      RECT 0.342 0.063 0.36 0.131 ;
      RECT 0.338 0.063 0.375 0.081 ;
      RECT 0.207 0.171 0.245 0.189 ;
      RECT 0.227 0.027 0.245 0.189 ;
      RECT 0.207 0.027 0.245 0.045 ;
      RECT 0.138 0.099 0.198 0.117 ;
      RECT 0.18 0.063 0.198 0.117 ;
      RECT 0.143 0.063 0.198 0.081 ;
      RECT 0.016 0.171 0.068 0.189 ;
      RECT 0.016 0.027 0.034 0.189 ;
      RECT 0.016 0.027 0.068 0.045 ;
      RECT 0.504 0.044 0.522 0.103 ;
    LAYER M2 ;
      RECT 0.45 0.135 0.61 0.153 ;
      RECT 0.016 0.063 0.527 0.081 ;
      RECT 0.222 0.135 0.414 0.153 ;
    LAYER V1 ;
      RECT 0.585 0.135 0.603 0.153 ;
      RECT 0.504 0.063 0.522 0.081 ;
      RECT 0.45 0.135 0.468 0.153 ;
      RECT 0.396 0.135 0.414 0.153 ;
      RECT 0.342 0.063 0.36 0.081 ;
      RECT 0.227 0.135 0.245 0.153 ;
      RECT 0.153 0.063 0.171 0.081 ;
      RECT 0.016 0.063 0.034 0.081 ;
  END
END DLLx3_ASAP7_6t_SL

MACRO FAxp33_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FAxp33_ASAP7_6t_SL 0 0 ;
  SIZE 0.756 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.756 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.756 0.009 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.063 0.649 0.081 ;
        RECT 0.612 0.063 0.63 0.125 ;
        RECT 0.389 0.099 0.431 0.117 ;
        RECT 0.413 0.058 0.431 0.117 ;
        RECT 0.018 0.063 0.078 0.081 ;
        RECT 0.018 0.063 0.036 0.13 ;
      LAYER M2 ;
        RECT 0.04 0.063 0.643 0.081 ;
      LAYER V1 ;
        RECT 0.045 0.063 0.063 0.081 ;
        RECT 0.413 0.063 0.431 0.081 ;
        RECT 0.618 0.063 0.636 0.081 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.686 0.171 0.738 0.189 ;
        RECT 0.72 0.088 0.738 0.189 ;
        RECT 0.31 0.171 0.365 0.189 ;
        RECT 0.31 0.094 0.328 0.189 ;
        RECT 0.18 0.135 0.328 0.153 ;
        RECT 0.18 0.094 0.198 0.153 ;
      LAYER M2 ;
        RECT 0.31 0.171 0.717 0.189 ;
      LAYER V1 ;
        RECT 0.315 0.171 0.333 0.189 ;
        RECT 0.693 0.171 0.711 0.189 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.543 0.099 0.586 0.117 ;
        RECT 0.543 0.079 0.561 0.125 ;
        RECT 0.45 0.092 0.468 0.145 ;
        RECT 0.237 0.099 0.292 0.117 ;
        RECT 0.274 0.063 0.292 0.117 ;
        RECT 0.237 0.063 0.292 0.081 ;
      LAYER M2 ;
        RECT 0.225 0.099 0.59 0.117 ;
      LAYER V1 ;
        RECT 0.252 0.099 0.27 0.117 ;
        RECT 0.45 0.099 0.468 0.117 ;
        RECT 0.564 0.099 0.582 0.117 ;
    END
  END CI
  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.501 0.072 0.519 0.135 ;
        RECT 0.486 0.117 0.504 0.172 ;
        RECT 0.124 0.038 0.208 0.056 ;
        RECT 0.14 0.135 0.158 0.176 ;
        RECT 0.124 0.038 0.142 0.153 ;
      LAYER M2 ;
        RECT 0.126 0.135 0.509 0.153 ;
      LAYER V1 ;
        RECT 0.134 0.135 0.152 0.153 ;
        RECT 0.486 0.135 0.504 0.153 ;
    END
  END CON
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.346 0.135 0.418 0.153 ;
        RECT 0.346 0.027 0.392 0.045 ;
        RECT 0.346 0.027 0.364 0.153 ;
      LAYER M2 ;
        RECT 0.363 0.027 0.649 0.045 ;
      LAYER V1 ;
        RECT 0.369 0.027 0.387 0.045 ;
    END
  END SN
  OBS
    LAYER M1 ;
      RECT 0.531 0.027 0.662 0.045 ;
      RECT 0.539 0.153 0.649 0.171 ;
      RECT 0.243 0.027 0.295 0.045 ;
      RECT 0.195 0.171 0.279 0.189 ;
      RECT 0.04 0.171 0.087 0.189 ;
      RECT 0.04 0.027 0.082 0.045 ;
    LAYER M2 ;
      RECT 0.04 0.027 0.284 0.045 ;
      RECT 0.04 0.171 0.231 0.189 ;
    LAYER V1 ;
      RECT 0.261 0.027 0.279 0.045 ;
      RECT 0.207 0.171 0.225 0.189 ;
      RECT 0.045 0.027 0.063 0.045 ;
      RECT 0.045 0.171 0.063 0.189 ;
  END
END FAxp33_ASAP7_6t_SL

MACRO FILLER_ASAP7_6t_SL
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN FILLER_ASAP7_6t_SL 0 0 ;
  SIZE 0.108 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.108 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.108 0.009 ;
    END
  END VSS
END FILLER_ASAP7_6t_SL

MACRO FILLERxp5_ASAP7_6t_SL
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN FILLERxp5_ASAP7_6t_SL 0 0 ;
  SIZE 0.054 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.054 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.054 0.009 ;
    END
  END VSS
END FILLERxp5_ASAP7_6t_SL

MACRO HAxp5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HAxp5_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.169 0.099 0.36 0.117 ;
        RECT 0.169 0.027 0.187 0.117 ;
        RECT 0.018 0.027 0.187 0.045 ;
        RECT 0.018 0.171 0.068 0.189 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.07 0.099 0.144 0.117 ;
        RECT 0.07 0.063 0.144 0.081 ;
        RECT 0.088 0.135 0.143 0.153 ;
        RECT 0.088 0.099 0.106 0.153 ;
        RECT 0.07 0.063 0.088 0.117 ;
    END
  END B
  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.176 0.135 0.414 0.153 ;
        RECT 0.396 0.063 0.414 0.153 ;
        RECT 0.212 0.063 0.414 0.081 ;
        RECT 0.099 0.171 0.194 0.189 ;
        RECT 0.176 0.135 0.194 0.189 ;
    END
  END CON
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.171 0.47 0.189 ;
        RECT 0.452 0.027 0.47 0.189 ;
        RECT 0.423 0.027 0.47 0.045 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.261 0.027 0.387 0.045 ;
  END
END HAxp5_ASAP7_6t_SL

MACRO HB1x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HB1x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.216 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.135 0.073 0.153 ;
        RECT 0.018 0.099 0.073 0.117 ;
        RECT 0.018 0.063 0.073 0.081 ;
        RECT 0.018 0.063 0.036 0.153 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.216 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.216 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.171 0.198 0.189 ;
        RECT 0.18 0.027 0.198 0.189 ;
        RECT 0.148 0.027 0.198 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.036 0.171 0.119 0.189 ;
      RECT 0.101 0.027 0.119 0.189 ;
      RECT 0.101 0.099 0.149 0.117 ;
      RECT 0.034 0.027 0.119 0.045 ;
  END
END HB1x1_ASAP7_6t_SL

MACRO HB2x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HB2x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.27 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.095 0.117 ;
        RECT 0.018 0.171 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.27 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.27 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.171 0.252 0.189 ;
        RECT 0.234 0.027 0.252 0.189 ;
        RECT 0.202 0.027 0.252 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.099 0.171 0.144 0.189 ;
      RECT 0.126 0.027 0.144 0.189 ;
      RECT 0.126 0.099 0.203 0.117 ;
      RECT 0.099 0.027 0.144 0.045 ;
  END
END HB2x1_ASAP7_6t_SL

MACRO HB3x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HB3x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.095 0.117 ;
        RECT 0.018 0.171 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.171 0.306 0.189 ;
        RECT 0.288 0.027 0.306 0.189 ;
        RECT 0.256 0.027 0.306 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.099 0.171 0.198 0.189 ;
      RECT 0.18 0.027 0.198 0.189 ;
      RECT 0.18 0.099 0.257 0.117 ;
      RECT 0.099 0.027 0.198 0.045 ;
  END
END HB3x1_ASAP7_6t_SL

MACRO HB4x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HB4x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.016 0.099 0.101 0.117 ;
        RECT 0.016 0.171 0.068 0.189 ;
        RECT 0.016 0.027 0.068 0.045 ;
        RECT 0.016 0.027 0.034 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.31 0.171 0.36 0.189 ;
        RECT 0.342 0.027 0.36 0.189 ;
        RECT 0.31 0.027 0.36 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.099 0.171 0.198 0.189 ;
      RECT 0.18 0.027 0.198 0.189 ;
      RECT 0.18 0.099 0.311 0.117 ;
      RECT 0.099 0.027 0.198 0.045 ;
  END
END HB4x1_ASAP7_6t_SL

MACRO ICGx10_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGx10_ASAP7_6t_SL 0 0 ;
  SIZE 1.674 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.93 0.135 0.986 0.153 ;
        RECT 0.968 0.11 0.986 0.153 ;
        RECT 0.612 0.135 0.76 0.153 ;
        RECT 0.742 0.11 0.76 0.153 ;
        RECT 0.649 0.027 0.706 0.045 ;
        RECT 0.612 0.063 0.667 0.081 ;
        RECT 0.649 0.027 0.667 0.081 ;
        RECT 0.612 0.063 0.63 0.153 ;
        RECT 0.396 0.113 0.414 0.172 ;
        RECT 0.23 0.135 0.267 0.153 ;
        RECT 0.234 0.085 0.252 0.153 ;
      LAYER M2 ;
        RECT 0.225 0.135 0.958 0.153 ;
      LAYER V1 ;
        RECT 0.234 0.135 0.252 0.153 ;
        RECT 0.396 0.135 0.414 0.153 ;
        RECT 0.668 0.135 0.686 0.153 ;
        RECT 0.94 0.135 0.958 0.153 ;
    END
  END CLK
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.098 0.09 0.116 ;
        RECT 0.018 0.171 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END ENA
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.098 0.171 1.631 0.189 ;
        RECT 1.611 0.027 1.631 0.189 ;
        RECT 1.101 0.027 1.631 0.045 ;
    END
  END GCLK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.135 0.144 0.153 ;
        RECT 0.126 0.063 0.144 0.153 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.674 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.674 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.685 0.171 1.062 0.189 ;
      RECT 1.044 0.135 1.062 0.189 ;
      RECT 1.044 0.135 1.116 0.153 ;
      RECT 1.098 0.063 1.116 0.153 ;
      RECT 1.048 0.063 1.116 0.081 ;
      RECT 1.048 0.027 1.066 0.081 ;
      RECT 0.747 0.027 1.066 0.045 ;
      RECT 0.787 0.099 0.852 0.117 ;
      RECT 0.657 0.099 0.715 0.117 ;
      RECT 0.697 0.063 0.715 0.117 ;
      RECT 0.787 0.063 0.805 0.117 ;
      RECT 0.697 0.063 0.805 0.081 ;
      RECT 0.559 0.171 0.639 0.189 ;
      RECT 0.559 0.027 0.577 0.189 ;
      RECT 0.559 0.027 0.603 0.045 ;
      RECT 0.472 0.171 0.534 0.189 ;
      RECT 0.516 0.027 0.534 0.189 ;
      RECT 0.396 0.07 0.444 0.088 ;
      RECT 0.426 0.027 0.444 0.088 ;
      RECT 0.426 0.027 0.534 0.045 ;
      RECT 0.256 0.171 0.36 0.189 ;
      RECT 0.342 0.027 0.36 0.189 ;
      RECT 0.305 0.027 0.36 0.045 ;
      RECT 0.288 0.063 0.306 0.126 ;
      RECT 0.274 0.063 0.316 0.081 ;
      RECT 0.099 0.171 0.198 0.189 ;
      RECT 0.18 0.027 0.198 0.189 ;
      RECT 0.099 0.027 0.198 0.045 ;
      RECT 1.019 0.099 1.073 0.117 ;
      RECT 0.462 0.07 0.48 0.126 ;
    LAYER M2 ;
      RECT 0.33 0.099 1.07 0.117 ;
      RECT 0.282 0.063 0.586 0.081 ;
    LAYER V1 ;
      RECT 1.042 0.099 1.06 0.117 ;
      RECT 0.668 0.099 0.686 0.117 ;
      RECT 0.559 0.063 0.577 0.081 ;
      RECT 0.462 0.099 0.48 0.117 ;
      RECT 0.342 0.099 0.36 0.117 ;
      RECT 0.288 0.063 0.306 0.081 ;
  END
END ICGx10_ASAP7_6t_SL

MACRO ICGx12_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGx12_ASAP7_6t_SL 0 0 ;
  SIZE 1.782 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.93 0.135 0.986 0.153 ;
        RECT 0.968 0.11 0.986 0.153 ;
        RECT 0.612 0.135 0.76 0.153 ;
        RECT 0.742 0.11 0.76 0.153 ;
        RECT 0.649 0.027 0.706 0.045 ;
        RECT 0.612 0.063 0.667 0.081 ;
        RECT 0.649 0.027 0.667 0.081 ;
        RECT 0.612 0.063 0.63 0.153 ;
        RECT 0.396 0.113 0.414 0.172 ;
        RECT 0.23 0.135 0.267 0.153 ;
        RECT 0.234 0.085 0.252 0.153 ;
      LAYER M2 ;
        RECT 0.225 0.135 0.958 0.153 ;
      LAYER V1 ;
        RECT 0.234 0.135 0.252 0.153 ;
        RECT 0.396 0.135 0.414 0.153 ;
        RECT 0.668 0.135 0.686 0.153 ;
        RECT 0.94 0.135 0.958 0.153 ;
    END
  END CLK
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.054 0.098 0.09 0.116 ;
        RECT 0.035 0.135 0.072 0.153 ;
        RECT 0.054 0.027 0.072 0.153 ;
        RECT 0.035 0.027 0.072 0.045 ;
    END
  END ENA
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.095 0.171 1.721 0.189 ;
        RECT 1.703 0.027 1.721 0.189 ;
        RECT 1.098 0.027 1.721 0.045 ;
    END
  END GCLK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.135 0.144 0.153 ;
        RECT 0.126 0.063 0.144 0.153 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.782 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.782 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.685 0.171 1.062 0.189 ;
      RECT 1.044 0.135 1.062 0.189 ;
      RECT 1.044 0.135 1.116 0.153 ;
      RECT 1.098 0.063 1.116 0.153 ;
      RECT 1.048 0.063 1.116 0.081 ;
      RECT 1.048 0.027 1.066 0.081 ;
      RECT 0.747 0.027 1.066 0.045 ;
      RECT 0.787 0.099 0.852 0.117 ;
      RECT 0.657 0.099 0.715 0.117 ;
      RECT 0.697 0.063 0.715 0.117 ;
      RECT 0.787 0.063 0.805 0.117 ;
      RECT 0.697 0.063 0.805 0.081 ;
      RECT 0.559 0.171 0.639 0.189 ;
      RECT 0.559 0.027 0.577 0.189 ;
      RECT 0.559 0.027 0.603 0.045 ;
      RECT 0.472 0.171 0.534 0.189 ;
      RECT 0.516 0.027 0.534 0.189 ;
      RECT 0.396 0.07 0.444 0.088 ;
      RECT 0.426 0.027 0.444 0.088 ;
      RECT 0.426 0.027 0.534 0.045 ;
      RECT 0.256 0.171 0.36 0.189 ;
      RECT 0.342 0.027 0.36 0.189 ;
      RECT 0.305 0.027 0.36 0.045 ;
      RECT 0.288 0.063 0.306 0.126 ;
      RECT 0.274 0.063 0.316 0.081 ;
      RECT 0.037 0.171 0.198 0.189 ;
      RECT 0.18 0.027 0.198 0.189 ;
      RECT 0.099 0.027 0.198 0.045 ;
      RECT 1.019 0.099 1.073 0.117 ;
      RECT 0.462 0.07 0.48 0.126 ;
    LAYER M2 ;
      RECT 0.33 0.099 1.07 0.117 ;
      RECT 0.282 0.063 0.586 0.081 ;
    LAYER V1 ;
      RECT 1.042 0.099 1.06 0.117 ;
      RECT 0.668 0.099 0.686 0.117 ;
      RECT 0.559 0.063 0.577 0.081 ;
      RECT 0.462 0.099 0.48 0.117 ;
      RECT 0.342 0.099 0.36 0.117 ;
      RECT 0.288 0.063 0.306 0.081 ;
  END
END ICGx12_ASAP7_6t_SL

MACRO ICGx1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGx1_ASAP7_6t_SL 0 0 ;
  SIZE 0.972 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.135 0.76 0.153 ;
        RECT 0.742 0.11 0.76 0.153 ;
        RECT 0.649 0.027 0.706 0.045 ;
        RECT 0.612 0.063 0.667 0.081 ;
        RECT 0.649 0.027 0.667 0.081 ;
        RECT 0.612 0.063 0.63 0.153 ;
        RECT 0.396 0.171 0.446 0.189 ;
        RECT 0.396 0.113 0.414 0.189 ;
        RECT 0.234 0.027 0.289 0.045 ;
        RECT 0.23 0.135 0.267 0.153 ;
        RECT 0.234 0.027 0.252 0.153 ;
      LAYER M2 ;
        RECT 0.225 0.135 0.692 0.153 ;
      LAYER V1 ;
        RECT 0.234 0.135 0.252 0.153 ;
        RECT 0.396 0.135 0.414 0.153 ;
        RECT 0.668 0.135 0.686 0.153 ;
    END
  END CLK
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.054 0.098 0.09 0.116 ;
        RECT 0.035 0.17 0.072 0.189 ;
        RECT 0.054 0.027 0.072 0.189 ;
        RECT 0.035 0.027 0.072 0.045 ;
    END
  END ENA
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.878 0.171 0.953 0.189 ;
        RECT 0.935 0.027 0.953 0.189 ;
        RECT 0.881 0.027 0.953 0.045 ;
    END
  END GCLK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.135 0.144 0.153 ;
        RECT 0.126 0.063 0.144 0.153 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.972 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.972 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.688 0.171 0.846 0.189 ;
      RECT 0.828 0.135 0.846 0.189 ;
      RECT 0.828 0.135 0.9 0.153 ;
      RECT 0.882 0.063 0.9 0.153 ;
      RECT 0.832 0.063 0.9 0.081 ;
      RECT 0.832 0.027 0.85 0.081 ;
      RECT 0.737 0.027 0.85 0.045 ;
      RECT 0.787 0.099 0.852 0.117 ;
      RECT 0.657 0.099 0.715 0.117 ;
      RECT 0.697 0.063 0.715 0.117 ;
      RECT 0.787 0.063 0.805 0.117 ;
      RECT 0.697 0.063 0.805 0.081 ;
      RECT 0.559 0.171 0.639 0.189 ;
      RECT 0.559 0.027 0.577 0.189 ;
      RECT 0.559 0.027 0.603 0.045 ;
      RECT 0.477 0.171 0.534 0.189 ;
      RECT 0.516 0.027 0.534 0.189 ;
      RECT 0.396 0.07 0.444 0.088 ;
      RECT 0.426 0.027 0.444 0.088 ;
      RECT 0.426 0.027 0.534 0.045 ;
      RECT 0.256 0.171 0.36 0.189 ;
      RECT 0.342 0.034 0.36 0.189 ;
      RECT 0.288 0.063 0.306 0.126 ;
      RECT 0.277 0.063 0.316 0.081 ;
      RECT 0.099 0.171 0.198 0.189 ;
      RECT 0.18 0.027 0.198 0.189 ;
      RECT 0.099 0.027 0.198 0.045 ;
      RECT 0.462 0.07 0.48 0.126 ;
    LAYER M2 ;
      RECT 0.33 0.099 0.692 0.117 ;
      RECT 0.282 0.063 0.586 0.081 ;
    LAYER V1 ;
      RECT 0.668 0.099 0.686 0.117 ;
      RECT 0.559 0.063 0.577 0.081 ;
      RECT 0.462 0.099 0.48 0.117 ;
      RECT 0.342 0.099 0.36 0.117 ;
      RECT 0.288 0.063 0.306 0.081 ;
  END
END ICGx1_ASAP7_6t_SL

MACRO ICGx2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGx2_ASAP7_6t_SL 0 0 ;
  SIZE 1.026 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.135 0.76 0.153 ;
        RECT 0.742 0.11 0.76 0.153 ;
        RECT 0.649 0.027 0.706 0.045 ;
        RECT 0.612 0.063 0.667 0.081 ;
        RECT 0.649 0.027 0.667 0.081 ;
        RECT 0.612 0.063 0.63 0.153 ;
        RECT 0.396 0.17 0.446 0.188 ;
        RECT 0.396 0.113 0.414 0.188 ;
        RECT 0.234 0.027 0.289 0.045 ;
        RECT 0.23 0.135 0.267 0.153 ;
        RECT 0.234 0.027 0.252 0.153 ;
      LAYER M2 ;
        RECT 0.225 0.135 0.692 0.153 ;
      LAYER V1 ;
        RECT 0.234 0.135 0.252 0.153 ;
        RECT 0.396 0.135 0.414 0.153 ;
        RECT 0.668 0.135 0.686 0.153 ;
    END
  END CLK
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.054 0.098 0.09 0.116 ;
        RECT 0.035 0.171 0.072 0.189 ;
        RECT 0.054 0.027 0.072 0.189 ;
        RECT 0.035 0.027 0.072 0.045 ;
    END
  END ENA
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.879 0.171 0.954 0.189 ;
        RECT 0.936 0.027 0.954 0.189 ;
        RECT 0.882 0.027 0.954 0.045 ;
    END
  END GCLK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.135 0.144 0.153 ;
        RECT 0.126 0.063 0.144 0.153 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.026 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.026 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.688 0.171 0.846 0.189 ;
      RECT 0.828 0.135 0.846 0.189 ;
      RECT 0.828 0.135 0.9 0.153 ;
      RECT 0.882 0.063 0.9 0.153 ;
      RECT 0.832 0.063 0.9 0.081 ;
      RECT 0.832 0.027 0.85 0.081 ;
      RECT 0.737 0.027 0.85 0.045 ;
      RECT 0.787 0.099 0.852 0.117 ;
      RECT 0.657 0.099 0.715 0.117 ;
      RECT 0.697 0.063 0.715 0.117 ;
      RECT 0.787 0.063 0.805 0.117 ;
      RECT 0.697 0.063 0.805 0.081 ;
      RECT 0.559 0.171 0.639 0.189 ;
      RECT 0.559 0.027 0.577 0.189 ;
      RECT 0.559 0.027 0.603 0.045 ;
      RECT 0.477 0.171 0.534 0.189 ;
      RECT 0.516 0.027 0.534 0.189 ;
      RECT 0.396 0.07 0.444 0.088 ;
      RECT 0.426 0.027 0.444 0.088 ;
      RECT 0.426 0.027 0.534 0.045 ;
      RECT 0.256 0.171 0.36 0.189 ;
      RECT 0.342 0.034 0.36 0.189 ;
      RECT 0.288 0.063 0.306 0.126 ;
      RECT 0.277 0.063 0.316 0.081 ;
      RECT 0.099 0.171 0.198 0.189 ;
      RECT 0.18 0.027 0.198 0.189 ;
      RECT 0.099 0.027 0.198 0.045 ;
      RECT 0.462 0.07 0.48 0.126 ;
    LAYER M2 ;
      RECT 0.33 0.099 0.692 0.117 ;
      RECT 0.282 0.063 0.586 0.081 ;
    LAYER V1 ;
      RECT 0.668 0.099 0.686 0.117 ;
      RECT 0.559 0.063 0.577 0.081 ;
      RECT 0.462 0.099 0.48 0.117 ;
      RECT 0.342 0.099 0.36 0.117 ;
      RECT 0.288 0.063 0.306 0.081 ;
  END
END ICGx2_ASAP7_6t_SL

MACRO ICGx3_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGx3_ASAP7_6t_SL 0 0 ;
  SIZE 1.08 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.135 0.76 0.153 ;
        RECT 0.742 0.11 0.76 0.153 ;
        RECT 0.649 0.027 0.706 0.045 ;
        RECT 0.612 0.063 0.667 0.081 ;
        RECT 0.649 0.027 0.667 0.081 ;
        RECT 0.612 0.063 0.63 0.153 ;
        RECT 0.396 0.171 0.446 0.189 ;
        RECT 0.396 0.113 0.414 0.189 ;
        RECT 0.234 0.027 0.289 0.045 ;
        RECT 0.23 0.135 0.267 0.153 ;
        RECT 0.234 0.027 0.252 0.153 ;
      LAYER M2 ;
        RECT 0.225 0.135 0.692 0.153 ;
      LAYER V1 ;
        RECT 0.234 0.135 0.252 0.153 ;
        RECT 0.396 0.135 0.414 0.153 ;
        RECT 0.668 0.135 0.686 0.153 ;
    END
  END CLK
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.054 0.098 0.09 0.116 ;
        RECT 0.035 0.171 0.072 0.189 ;
        RECT 0.054 0.027 0.072 0.189 ;
        RECT 0.035 0.027 0.072 0.045 ;
    END
  END ENA
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.879 0.171 1.041 0.189 ;
        RECT 0.882 0.027 1.041 0.045 ;
        RECT 0.936 0.027 0.954 0.189 ;
    END
  END GCLK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.135 0.144 0.153 ;
        RECT 0.126 0.063 0.144 0.153 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.08 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.08 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.688 0.171 0.846 0.189 ;
      RECT 0.828 0.135 0.846 0.189 ;
      RECT 0.828 0.135 0.9 0.153 ;
      RECT 0.882 0.063 0.9 0.153 ;
      RECT 0.832 0.063 0.9 0.081 ;
      RECT 0.832 0.027 0.85 0.081 ;
      RECT 0.737 0.027 0.85 0.045 ;
      RECT 0.787 0.099 0.852 0.117 ;
      RECT 0.657 0.099 0.715 0.117 ;
      RECT 0.697 0.063 0.715 0.117 ;
      RECT 0.787 0.063 0.805 0.117 ;
      RECT 0.697 0.063 0.805 0.081 ;
      RECT 0.559 0.171 0.639 0.189 ;
      RECT 0.559 0.027 0.577 0.189 ;
      RECT 0.559 0.027 0.603 0.045 ;
      RECT 0.477 0.171 0.534 0.189 ;
      RECT 0.516 0.027 0.534 0.189 ;
      RECT 0.396 0.07 0.444 0.088 ;
      RECT 0.426 0.027 0.444 0.088 ;
      RECT 0.426 0.027 0.534 0.045 ;
      RECT 0.256 0.171 0.36 0.189 ;
      RECT 0.342 0.034 0.36 0.189 ;
      RECT 0.288 0.063 0.306 0.126 ;
      RECT 0.277 0.063 0.316 0.081 ;
      RECT 0.099 0.171 0.198 0.189 ;
      RECT 0.18 0.027 0.198 0.189 ;
      RECT 0.099 0.027 0.198 0.045 ;
      RECT 0.462 0.07 0.48 0.126 ;
    LAYER M2 ;
      RECT 0.33 0.099 0.692 0.117 ;
      RECT 0.282 0.063 0.586 0.081 ;
    LAYER V1 ;
      RECT 0.668 0.099 0.686 0.117 ;
      RECT 0.559 0.063 0.577 0.081 ;
      RECT 0.462 0.099 0.48 0.117 ;
      RECT 0.342 0.099 0.36 0.117 ;
      RECT 0.288 0.063 0.306 0.081 ;
  END
END ICGx3_ASAP7_6t_SL

MACRO ICGx4_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGx4_ASAP7_6t_SL 0 0 ;
  SIZE 1.35 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.93 0.135 0.986 0.153 ;
        RECT 0.968 0.11 0.986 0.153 ;
        RECT 0.612 0.135 0.76 0.153 ;
        RECT 0.742 0.11 0.76 0.153 ;
        RECT 0.649 0.027 0.706 0.045 ;
        RECT 0.612 0.063 0.667 0.081 ;
        RECT 0.649 0.027 0.667 0.081 ;
        RECT 0.612 0.063 0.63 0.153 ;
        RECT 0.396 0.171 0.446 0.189 ;
        RECT 0.396 0.113 0.414 0.189 ;
        RECT 0.233 0.027 0.292 0.045 ;
        RECT 0.23 0.135 0.267 0.153 ;
        RECT 0.234 0.027 0.252 0.153 ;
      LAYER M2 ;
        RECT 0.225 0.135 0.958 0.153 ;
      LAYER V1 ;
        RECT 0.234 0.135 0.252 0.153 ;
        RECT 0.396 0.135 0.414 0.153 ;
        RECT 0.668 0.135 0.686 0.153 ;
        RECT 0.94 0.135 0.958 0.153 ;
    END
  END CLK
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.054 0.098 0.09 0.116 ;
        RECT 0.035 0.171 0.072 0.189 ;
        RECT 0.054 0.027 0.072 0.189 ;
        RECT 0.035 0.027 0.072 0.045 ;
    END
  END ENA
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.095 0.171 1.294 0.189 ;
        RECT 1.276 0.027 1.294 0.189 ;
        RECT 1.098 0.027 1.294 0.045 ;
    END
  END GCLK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.135 0.144 0.153 ;
        RECT 0.126 0.063 0.144 0.153 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.35 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.35 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.685 0.171 1.062 0.189 ;
      RECT 1.044 0.135 1.062 0.189 ;
      RECT 1.044 0.135 1.116 0.153 ;
      RECT 1.098 0.063 1.116 0.153 ;
      RECT 1.048 0.063 1.116 0.081 ;
      RECT 1.048 0.027 1.066 0.081 ;
      RECT 0.747 0.027 1.066 0.045 ;
      RECT 0.787 0.099 0.852 0.117 ;
      RECT 0.657 0.099 0.715 0.117 ;
      RECT 0.697 0.063 0.715 0.117 ;
      RECT 0.787 0.063 0.805 0.117 ;
      RECT 0.697 0.063 0.805 0.081 ;
      RECT 0.559 0.171 0.639 0.189 ;
      RECT 0.559 0.027 0.577 0.189 ;
      RECT 0.559 0.027 0.603 0.045 ;
      RECT 0.477 0.171 0.534 0.189 ;
      RECT 0.516 0.027 0.534 0.189 ;
      RECT 0.396 0.07 0.444 0.088 ;
      RECT 0.426 0.027 0.444 0.088 ;
      RECT 0.426 0.027 0.534 0.045 ;
      RECT 0.256 0.171 0.36 0.189 ;
      RECT 0.342 0.034 0.36 0.189 ;
      RECT 0.288 0.063 0.306 0.126 ;
      RECT 0.277 0.063 0.316 0.081 ;
      RECT 0.099 0.171 0.198 0.189 ;
      RECT 0.18 0.027 0.198 0.189 ;
      RECT 0.099 0.027 0.198 0.045 ;
      RECT 1.019 0.099 1.073 0.117 ;
      RECT 0.462 0.07 0.48 0.126 ;
    LAYER M2 ;
      RECT 0.33 0.099 1.07 0.117 ;
      RECT 0.282 0.063 0.586 0.081 ;
    LAYER V1 ;
      RECT 1.042 0.099 1.06 0.117 ;
      RECT 0.668 0.099 0.686 0.117 ;
      RECT 0.559 0.063 0.577 0.081 ;
      RECT 0.462 0.099 0.48 0.117 ;
      RECT 0.342 0.099 0.36 0.117 ;
      RECT 0.288 0.063 0.306 0.081 ;
  END
END ICGx4_ASAP7_6t_SL

MACRO ICGx5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGx5_ASAP7_6t_SL 0 0 ;
  SIZE 1.404 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.93 0.135 0.986 0.153 ;
        RECT 0.968 0.11 0.986 0.153 ;
        RECT 0.612 0.135 0.76 0.153 ;
        RECT 0.742 0.11 0.76 0.153 ;
        RECT 0.649 0.027 0.706 0.045 ;
        RECT 0.612 0.063 0.667 0.081 ;
        RECT 0.649 0.027 0.667 0.081 ;
        RECT 0.612 0.063 0.63 0.153 ;
        RECT 0.396 0.171 0.446 0.189 ;
        RECT 0.396 0.113 0.414 0.189 ;
        RECT 0.234 0.027 0.289 0.045 ;
        RECT 0.23 0.135 0.267 0.153 ;
        RECT 0.234 0.027 0.252 0.153 ;
      LAYER M2 ;
        RECT 0.225 0.135 0.958 0.153 ;
      LAYER V1 ;
        RECT 0.234 0.135 0.252 0.153 ;
        RECT 0.396 0.135 0.414 0.153 ;
        RECT 0.668 0.135 0.686 0.153 ;
        RECT 0.94 0.135 0.958 0.153 ;
    END
  END CLK
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.054 0.098 0.09 0.116 ;
        RECT 0.035 0.17 0.072 0.189 ;
        RECT 0.054 0.027 0.072 0.189 ;
        RECT 0.035 0.027 0.072 0.045 ;
    END
  END ENA
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.095 0.171 1.382 0.189 ;
        RECT 1.364 0.027 1.382 0.189 ;
        RECT 1.098 0.027 1.382 0.045 ;
    END
  END GCLK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.135 0.144 0.153 ;
        RECT 0.126 0.063 0.144 0.153 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.404 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.404 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.685 0.171 1.062 0.189 ;
      RECT 1.044 0.135 1.062 0.189 ;
      RECT 1.044 0.135 1.116 0.153 ;
      RECT 1.098 0.063 1.116 0.153 ;
      RECT 1.048 0.063 1.116 0.081 ;
      RECT 1.048 0.027 1.066 0.081 ;
      RECT 0.747 0.027 1.066 0.045 ;
      RECT 0.787 0.099 0.852 0.117 ;
      RECT 0.657 0.099 0.715 0.117 ;
      RECT 0.697 0.063 0.715 0.117 ;
      RECT 0.787 0.063 0.805 0.117 ;
      RECT 0.697 0.063 0.805 0.081 ;
      RECT 0.559 0.171 0.639 0.189 ;
      RECT 0.559 0.027 0.577 0.189 ;
      RECT 0.559 0.027 0.603 0.045 ;
      RECT 0.477 0.171 0.534 0.189 ;
      RECT 0.516 0.027 0.534 0.189 ;
      RECT 0.396 0.07 0.444 0.088 ;
      RECT 0.426 0.027 0.444 0.088 ;
      RECT 0.426 0.027 0.534 0.045 ;
      RECT 0.256 0.171 0.36 0.189 ;
      RECT 0.342 0.034 0.36 0.189 ;
      RECT 0.288 0.063 0.306 0.126 ;
      RECT 0.277 0.063 0.316 0.081 ;
      RECT 0.099 0.171 0.198 0.189 ;
      RECT 0.18 0.027 0.198 0.189 ;
      RECT 0.099 0.027 0.198 0.045 ;
      RECT 1.019 0.099 1.073 0.117 ;
      RECT 0.462 0.07 0.48 0.126 ;
    LAYER M2 ;
      RECT 0.33 0.099 1.07 0.117 ;
      RECT 0.282 0.063 0.586 0.081 ;
    LAYER V1 ;
      RECT 1.042 0.099 1.06 0.117 ;
      RECT 0.668 0.099 0.686 0.117 ;
      RECT 0.559 0.063 0.577 0.081 ;
      RECT 0.462 0.099 0.48 0.117 ;
      RECT 0.342 0.099 0.36 0.117 ;
      RECT 0.288 0.063 0.306 0.081 ;
  END
END ICGx5_ASAP7_6t_SL

MACRO ICGx8_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGx8_ASAP7_6t_SL 0 0 ;
  SIZE 1.566 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.93 0.135 0.986 0.153 ;
        RECT 0.968 0.11 0.986 0.153 ;
        RECT 0.612 0.135 0.76 0.153 ;
        RECT 0.742 0.11 0.76 0.153 ;
        RECT 0.649 0.027 0.716 0.045 ;
        RECT 0.612 0.063 0.667 0.081 ;
        RECT 0.649 0.027 0.667 0.081 ;
        RECT 0.612 0.063 0.63 0.153 ;
        RECT 0.396 0.113 0.414 0.172 ;
        RECT 0.23 0.135 0.267 0.153 ;
        RECT 0.234 0.085 0.252 0.153 ;
      LAYER M2 ;
        RECT 0.225 0.135 0.958 0.153 ;
      LAYER V1 ;
        RECT 0.234 0.135 0.252 0.153 ;
        RECT 0.396 0.135 0.414 0.153 ;
        RECT 0.668 0.135 0.686 0.153 ;
        RECT 0.94 0.135 0.958 0.153 ;
    END
  END CLK
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.098 0.095 0.116 ;
        RECT 0.018 0.171 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END ENA
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.12 0.171 1.508 0.189 ;
        RECT 1.49 0.027 1.508 0.189 ;
        RECT 1.12 0.027 1.508 0.045 ;
    END
  END GCLK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.135 0.144 0.153 ;
        RECT 0.126 0.063 0.144 0.153 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.566 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.566 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.685 0.171 1.062 0.189 ;
      RECT 1.044 0.135 1.062 0.189 ;
      RECT 1.044 0.135 1.109 0.153 ;
      RECT 1.091 0.063 1.109 0.153 ;
      RECT 1.091 0.1 1.364 0.118 ;
      RECT 1.048 0.063 1.109 0.081 ;
      RECT 1.048 0.027 1.066 0.081 ;
      RECT 0.747 0.027 1.066 0.045 ;
      RECT 0.787 0.099 0.852 0.117 ;
      RECT 0.657 0.099 0.715 0.117 ;
      RECT 0.697 0.063 0.715 0.117 ;
      RECT 0.787 0.063 0.805 0.117 ;
      RECT 0.697 0.063 0.805 0.081 ;
      RECT 0.552 0.171 0.603 0.189 ;
      RECT 0.552 0.027 0.57 0.189 ;
      RECT 0.552 0.027 0.603 0.045 ;
      RECT 0.472 0.171 0.534 0.189 ;
      RECT 0.516 0.027 0.534 0.189 ;
      RECT 0.396 0.07 0.444 0.088 ;
      RECT 0.426 0.027 0.444 0.088 ;
      RECT 0.426 0.027 0.534 0.045 ;
      RECT 0.256 0.171 0.36 0.189 ;
      RECT 0.342 0.027 0.36 0.189 ;
      RECT 0.305 0.027 0.36 0.045 ;
      RECT 0.288 0.063 0.306 0.126 ;
      RECT 0.274 0.063 0.316 0.081 ;
      RECT 0.099 0.171 0.198 0.189 ;
      RECT 0.18 0.027 0.198 0.189 ;
      RECT 0.099 0.027 0.198 0.045 ;
      RECT 1.019 0.099 1.066 0.117 ;
      RECT 0.462 0.07 0.48 0.126 ;
    LAYER M2 ;
      RECT 0.33 0.099 1.07 0.117 ;
      RECT 0.283 0.063 0.575 0.081 ;
    LAYER V1 ;
      RECT 1.042 0.099 1.06 0.117 ;
      RECT 0.668 0.099 0.686 0.117 ;
      RECT 0.552 0.063 0.57 0.081 ;
      RECT 0.462 0.099 0.48 0.117 ;
      RECT 0.342 0.099 0.36 0.117 ;
      RECT 0.288 0.063 0.306 0.081 ;
  END
END ICGx8_ASAP7_6t_SL

MACRO INVx11_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx11_ASAP7_6t_SL 0 0 ;
  SIZE 0.702 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.078 0.117 ;
        RECT 0.018 0.152 0.069 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.702 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.702 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.684 0.189 ;
        RECT 0.666 0.027 0.684 0.189 ;
        RECT 0.094 0.027 0.684 0.045 ;
    END
  END Y
END INVx11_ASAP7_6t_SL

MACRO INVx13_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx13_ASAP7_6t_SL 0 0 ;
  SIZE 0.81 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.078 0.117 ;
        RECT 0.018 0.171 0.055 0.189 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.81 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.81 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.792 0.189 ;
        RECT 0.774 0.027 0.792 0.189 ;
        RECT 0.094 0.027 0.792 0.045 ;
    END
  END Y
END INVx13_ASAP7_6t_SL

MACRO INVx1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx1_ASAP7_6t_SL 0 0 ;
  SIZE 0.162 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.078 0.117 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.162 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.162 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.144 0.189 ;
        RECT 0.126 0.027 0.144 0.189 ;
        RECT 0.094 0.027 0.144 0.045 ;
    END
  END Y
END INVx1_ASAP7_6t_SL

MACRO INVx2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx2_ASAP7_6t_SL 0 0 ;
  SIZE 0.216 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.216 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.216 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.198 0.189 ;
        RECT 0.18 0.027 0.198 0.189 ;
        RECT 0.094 0.027 0.198 0.045 ;
    END
  END Y
END INVx2_ASAP7_6t_SL

MACRO INVx3_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx3_ASAP7_6t_SL 0 0 ;
  SIZE 0.27 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.078 0.117 ;
        RECT 0.018 0.152 0.069 0.189 ;
        RECT 0.018 0.027 0.069 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.27 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.27 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.252 0.189 ;
        RECT 0.234 0.027 0.252 0.189 ;
        RECT 0.094 0.027 0.252 0.045 ;
    END
  END Y
END INVx3_ASAP7_6t_SL

MACRO INVx4_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx4_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.078 0.117 ;
        RECT 0.018 0.171 0.055 0.189 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.306 0.189 ;
        RECT 0.288 0.027 0.306 0.189 ;
        RECT 0.094 0.027 0.306 0.045 ;
    END
  END Y
END INVx4_ASAP7_6t_SL

MACRO INVx5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx5_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.095 0.117 ;
        RECT 0.018 0.171 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.171 0.36 0.189 ;
        RECT 0.342 0.027 0.36 0.189 ;
        RECT 0.099 0.027 0.36 0.045 ;
    END
  END Y
END INVx5_ASAP7_6t_SL

MACRO INVx6_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx6_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.078 0.117 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.414 0.189 ;
        RECT 0.396 0.027 0.414 0.189 ;
        RECT 0.094 0.027 0.414 0.045 ;
    END
  END Y
END INVx6_ASAP7_6t_SL

MACRO INVx8_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx8_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.078 0.117 ;
        RECT 0.018 0.152 0.069 0.189 ;
        RECT 0.018 0.027 0.069 0.072 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.522 0.189 ;
        RECT 0.504 0.027 0.522 0.189 ;
        RECT 0.094 0.027 0.522 0.045 ;
    END
  END Y
END INVx8_ASAP7_6t_SL

MACRO INVxp5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVxp5_ASAP7_6t_SL 0 0 ;
  SIZE 0.162 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.078 0.117 ;
        RECT 0.018 0.171 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.162 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.162 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.171 0.144 0.189 ;
        RECT 0.126 0.027 0.144 0.189 ;
        RECT 0.099 0.027 0.144 0.045 ;
    END
  END Y
END INVxp5_ASAP7_6t_SL

MACRO MAJIxp5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MAJIxp5_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.054 0.099 0.178 0.117 ;
        RECT 0.035 0.171 0.072 0.189 ;
        RECT 0.054 0.099 0.072 0.189 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.291 0.135 0.402 0.153 ;
        RECT 0.291 0.063 0.351 0.081 ;
        RECT 0.291 0.063 0.309 0.153 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.171 0.403 0.189 ;
        RECT 0.145 0.027 0.333 0.045 ;
        RECT 0.255 0.027 0.273 0.189 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.027 0.393 0.045 ;
      LAYER M1 ;
        RECT 0.386 0.099 0.423 0.117 ;
        RECT 0.405 0.027 0.423 0.117 ;
        RECT 0.364 0.027 0.423 0.045 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.123 ;
      LAYER V1 ;
        RECT 0.045 0.027 0.063 0.045 ;
        RECT 0.369 0.027 0.387 0.045 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.093 0.063 0.23 0.081 ;
      RECT 0.099 0.135 0.23 0.153 ;
  END
END MAJIxp5_ASAP7_6t_SL

MACRO MAJx1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MAJx1_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.127 0.135 0.182 0.153 ;
        RECT 0.164 0.063 0.182 0.153 ;
        RECT 0.127 0.063 0.182 0.081 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.171 0.357 0.189 ;
        RECT 0.339 0.09 0.357 0.189 ;
        RECT 0.018 0.063 0.056 0.081 ;
        RECT 0.018 0.063 0.036 0.189 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.135 0.252 0.153 ;
        RECT 0.234 0.063 0.252 0.153 ;
        RECT 0.207 0.063 0.252 0.081 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.418 0.171 0.468 0.189 ;
        RECT 0.45 0.027 0.468 0.189 ;
        RECT 0.418 0.027 0.468 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.28 0.135 0.321 0.153 ;
      RECT 0.303 0.027 0.321 0.153 ;
      RECT 0.061 0.135 0.102 0.153 ;
      RECT 0.084 0.027 0.102 0.153 ;
      RECT 0.375 0.099 0.412 0.117 ;
      RECT 0.375 0.027 0.393 0.117 ;
      RECT 0.028 0.027 0.393 0.045 ;
  END
END MAJx1_ASAP7_6t_SL

MACRO MAJx2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MAJx2_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.127 0.135 0.182 0.153 ;
        RECT 0.164 0.063 0.182 0.153 ;
        RECT 0.127 0.063 0.182 0.081 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.171 0.357 0.189 ;
        RECT 0.339 0.09 0.357 0.189 ;
        RECT 0.018 0.063 0.056 0.081 ;
        RECT 0.018 0.063 0.036 0.189 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.135 0.252 0.153 ;
        RECT 0.234 0.063 0.252 0.153 ;
        RECT 0.207 0.063 0.252 0.081 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.418 0.171 0.468 0.189 ;
        RECT 0.45 0.027 0.468 0.189 ;
        RECT 0.418 0.027 0.468 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.28 0.135 0.321 0.153 ;
      RECT 0.303 0.027 0.321 0.153 ;
      RECT 0.061 0.135 0.102 0.153 ;
      RECT 0.084 0.027 0.102 0.153 ;
      RECT 0.375 0.099 0.412 0.117 ;
      RECT 0.375 0.027 0.393 0.117 ;
      RECT 0.028 0.027 0.393 0.045 ;
  END
END MAJx2_ASAP7_6t_SL

MACRO MAJx3_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MAJx3_ASAP7_6t_SL 0 0 ;
  SIZE 0.594 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.127 0.135 0.182 0.153 ;
        RECT 0.164 0.063 0.182 0.153 ;
        RECT 0.127 0.063 0.182 0.081 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.171 0.357 0.189 ;
        RECT 0.339 0.09 0.357 0.189 ;
        RECT 0.018 0.063 0.056 0.081 ;
        RECT 0.018 0.063 0.036 0.189 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.135 0.252 0.153 ;
        RECT 0.234 0.063 0.252 0.153 ;
        RECT 0.207 0.063 0.252 0.081 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.594 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.418 0.171 0.555 0.189 ;
        RECT 0.418 0.027 0.555 0.045 ;
        RECT 0.45 0.027 0.468 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.28 0.135 0.321 0.153 ;
      RECT 0.303 0.027 0.321 0.153 ;
      RECT 0.061 0.135 0.102 0.153 ;
      RECT 0.084 0.027 0.102 0.153 ;
      RECT 0.375 0.099 0.412 0.117 ;
      RECT 0.375 0.027 0.393 0.117 ;
      RECT 0.028 0.027 0.393 0.045 ;
  END
END MAJx3_ASAP7_6t_SL

MACRO NAND2x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.084 0.117 ;
        RECT 0.018 0.063 0.073 0.081 ;
        RECT 0.018 0.171 0.068 0.189 ;
        RECT 0.018 0.063 0.036 0.189 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.115 0.099 0.23 0.117 ;
        RECT 0.115 0.135 0.17 0.153 ;
        RECT 0.115 0.063 0.17 0.081 ;
        RECT 0.115 0.063 0.133 0.153 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.171 0.311 0.189 ;
        RECT 0.293 0.063 0.311 0.189 ;
        RECT 0.202 0.063 0.311 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.027 0.284 0.045 ;
  END
END NAND2x1_ASAP7_6t_SL

MACRO NAND2x1p5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2x1p5_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.084 0.117 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.117 0.135 0.338 0.153 ;
        RECT 0.117 0.099 0.284 0.117 ;
        RECT 0.117 0.063 0.172 0.081 ;
        RECT 0.117 0.063 0.135 0.153 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.414 0.189 ;
        RECT 0.396 0.027 0.414 0.189 ;
        RECT 0.261 0.027 0.414 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.207 0.063 0.338 0.081 ;
      RECT 0.094 0.027 0.23 0.045 ;
  END
END NAND2x1p5_ASAP7_6t_SL

MACRO NAND2x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.135 0.297 0.153 ;
        RECT 0.279 0.099 0.297 0.153 ;
        RECT 0.242 0.099 0.297 0.117 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.413 0.135 0.468 0.153 ;
        RECT 0.45 0.099 0.468 0.153 ;
        RECT 0.322 0.099 0.468 0.117 ;
        RECT 0.322 0.063 0.34 0.117 ;
        RECT 0.182 0.063 0.34 0.081 ;
        RECT 0.072 0.099 0.2 0.117 ;
        RECT 0.182 0.063 0.2 0.117 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.171 0.522 0.189 ;
        RECT 0.504 0.063 0.522 0.189 ;
        RECT 0.418 0.063 0.522 0.081 ;
        RECT 0.018 0.063 0.122 0.081 ;
        RECT 0.018 0.063 0.036 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.027 0.5 0.045 ;
  END
END NAND2x2_ASAP7_6t_SL

MACRO NAND2xp5R_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2xp5R_ASAP7_6t_SL 0 0 ;
  SIZE 0.216 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.031 0.171 0.068 0.189 ;
        RECT 0.05 0.027 0.068 0.189 ;
        RECT 0.031 0.027 0.068 0.045 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.105 0.135 0.16 0.153 ;
        RECT 0.105 0.099 0.16 0.117 ;
        RECT 0.105 0.027 0.123 0.153 ;
        RECT 0.086 0.027 0.123 0.064 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.216 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.216 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.207 0.189 ;
        RECT 0.189 0.027 0.207 0.189 ;
        RECT 0.148 0.027 0.207 0.045 ;
    END
  END Y
END NAND2xp5R_ASAP7_6t_SL

MACRO NAND2xp5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2xp5_ASAP7_6t_SL 0 0 ;
  SIZE 0.216 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.171 0.068 0.189 ;
        RECT 0.017 0.027 0.068 0.064 ;
        RECT 0.017 0.027 0.035 0.189 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.089 0.099 0.144 0.117 ;
        RECT 0.089 0.027 0.126 0.153 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.216 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.216 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.171 0.198 0.189 ;
        RECT 0.18 0.027 0.198 0.189 ;
        RECT 0.148 0.027 0.198 0.064 ;
    END
  END Y
END NAND2xp5_ASAP7_6t_SL

MACRO NAND3x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.594 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.371 0.135 0.453 0.153 ;
        RECT 0.371 0.099 0.452 0.117 ;
        RECT 0.371 0.099 0.389 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.128 0.099 0.338 0.117 ;
        RECT 0.128 0.063 0.197 0.081 ;
        RECT 0.128 0.148 0.177 0.189 ;
        RECT 0.128 0.063 0.146 0.189 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.084 0.117 ;
        RECT 0.018 0.171 0.08 0.189 ;
        RECT 0.018 0.027 0.068 0.07 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.594 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.171 0.576 0.189 ;
        RECT 0.558 0.027 0.576 0.189 ;
        RECT 0.418 0.027 0.576 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.256 0.063 0.5 0.081 ;
      RECT 0.094 0.027 0.338 0.045 ;
  END
END NAND3x1_ASAP7_6t_SL

MACRO NAND3x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3x2_ASAP7_6t_SL 0 0 ;
  SIZE 1.08 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.153 0.135 1.001 0.153 ;
        RECT 0.983 0.099 1.001 0.153 ;
        RECT 0.891 0.099 1.001 0.117 ;
        RECT 0.153 0.099 0.171 0.153 ;
        RECT 0.094 0.099 0.171 0.117 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.519 0.063 0.579 0.081 ;
        RECT 0.519 0.099 0.575 0.117 ;
        RECT 0.519 0.063 0.537 0.117 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.08 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.08 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.171 1.062 0.189 ;
        RECT 1.044 0.027 1.062 0.189 ;
        RECT 0.904 0.027 1.062 0.045 ;
        RECT 0.018 0.027 0.176 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.31 0.099 0.752 0.117 ;
      LAYER M1 ;
        RECT 0.651 0.099 0.752 0.117 ;
        RECT 0.651 0.063 0.711 0.081 ;
        RECT 0.651 0.063 0.669 0.117 ;
        RECT 0.31 0.099 0.429 0.117 ;
        RECT 0.411 0.063 0.429 0.117 ;
        RECT 0.369 0.063 0.429 0.081 ;
      LAYER V1 ;
        RECT 0.315 0.099 0.333 0.117 ;
        RECT 0.729 0.099 0.747 0.117 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.742 0.063 0.986 0.081 ;
      RECT 0.256 0.027 0.824 0.045 ;
      RECT 0.094 0.063 0.338 0.081 ;
  END
END NAND3x2_ASAP7_6t_SL

MACRO NAND3xp33R_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3xp33R_ASAP7_6t_SL 0 0 ;
  SIZE 0.27 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.086 0.135 0.123 0.153 ;
        RECT 0.086 0.027 0.123 0.064 ;
        RECT 0.086 0.027 0.104 0.153 ;
        RECT 0.068 0.1 0.104 0.118 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.135 0.185 0.153 ;
        RECT 0.147 0.027 0.184 0.064 ;
        RECT 0.148 0.027 0.166 0.153 ;
        RECT 0.129 0.096 0.166 0.114 ;
        RECT 0.147 0.027 0.166 0.114 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.171 0.252 0.189 ;
        RECT 0.234 0.027 0.252 0.189 ;
        RECT 0.202 0.027 0.252 0.064 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.27 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.27 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.024 0.171 0.171 0.189 ;
        RECT 0.024 0.027 0.068 0.064 ;
        RECT 0.024 0.027 0.042 0.189 ;
    END
  END Y
END NAND3xp33R_ASAP7_6t_SL

MACRO NAND3xp33_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3xp33_ASAP7_6t_SL 0 0 ;
  SIZE 0.27 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.054 0.135 0.095 0.153 ;
        RECT 0.054 0.063 0.095 0.081 ;
        RECT 0.054 0.063 0.072 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.027 0.176 0.064 ;
        RECT 0.126 0.135 0.163 0.153 ;
        RECT 0.126 0.027 0.144 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.151 0.252 0.189 ;
        RECT 0.234 0.027 0.252 0.189 ;
        RECT 0.178 0.099 0.252 0.117 ;
        RECT 0.203 0.027 0.252 0.064 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.27 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.27 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.171 0.176 0.189 ;
        RECT 0.018 0.027 0.073 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END Y
END NAND3xp33_ASAP7_6t_SL

MACRO NAND4xp25R_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4xp25R_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.116 0.279 0.153 ;
        RECT 0.261 0.063 0.279 0.153 ;
        RECT 0.234 0.063 0.279 0.081 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.162 0.135 0.217 0.153 ;
        RECT 0.162 0.099 0.217 0.117 ;
        RECT 0.162 0.027 0.216 0.045 ;
        RECT 0.162 0.027 0.18 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.135 0.144 0.153 ;
        RECT 0.126 0.027 0.144 0.153 ;
        RECT 0.094 0.027 0.144 0.064 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.019 0.135 0.074 0.153 ;
        RECT 0.019 0.099 0.074 0.117 ;
        RECT 0.019 0.027 0.068 0.064 ;
        RECT 0.019 0.027 0.037 0.153 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.04 0.171 0.315 0.189 ;
        RECT 0.297 0.027 0.315 0.189 ;
        RECT 0.256 0.027 0.315 0.045 ;
    END
  END Y
END NAND4xp25R_ASAP7_6t_SL

MACRO NAND4xp25_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4xp25_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.225 0.135 0.27 0.153 ;
        RECT 0.252 0.09 0.27 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.162 0.027 0.23 0.064 ;
        RECT 0.162 0.099 0.207 0.117 ;
        RECT 0.162 0.027 0.18 0.146 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.135 0.144 0.153 ;
        RECT 0.126 0.027 0.144 0.153 ;
        RECT 0.09 0.027 0.144 0.07 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.135 0.073 0.153 ;
        RECT 0.018 0.099 0.073 0.117 ;
        RECT 0.018 0.027 0.068 0.07 ;
        RECT 0.018 0.027 0.036 0.153 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.04 0.171 0.306 0.189 ;
        RECT 0.288 0.027 0.306 0.189 ;
        RECT 0.256 0.027 0.306 0.045 ;
    END
  END Y
END NAND4xp25_ASAP7_6t_SL

MACRO NAND4xp75_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4xp75_ASAP7_6t_SL 0 0 ;
  SIZE 0.756 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.627 0.135 0.683 0.153 ;
        RECT 0.665 0.099 0.683 0.153 ;
        RECT 0.628 0.099 0.683 0.117 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.472 0.135 0.55 0.153 ;
        RECT 0.531 0.099 0.549 0.153 ;
        RECT 0.472 0.099 0.549 0.117 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.135 0.334 0.153 ;
        RECT 0.316 0.099 0.334 0.153 ;
        RECT 0.256 0.099 0.334 0.117 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.176 0.117 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.756 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.756 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.738 0.189 ;
        RECT 0.72 0.027 0.738 0.189 ;
        RECT 0.58 0.027 0.738 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.418 0.063 0.662 0.081 ;
      RECT 0.256 0.027 0.5 0.045 ;
      RECT 0.094 0.063 0.338 0.081 ;
  END
END NAND4xp75_ASAP7_6t_SL

MACRO NAND5xp2R_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND5xp2R_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.135 0.082 0.153 ;
        RECT 0.045 0.07 0.063 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.125 0.027 0.143 0.116 ;
        RECT 0.094 0.027 0.143 0.064 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.027 0.23 0.064 ;
        RECT 0.18 0.135 0.217 0.153 ;
        RECT 0.18 0.027 0.198 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.255 0.116 0.292 0.153 ;
        RECT 0.255 0.027 0.292 0.064 ;
        RECT 0.232 0.098 0.273 0.116 ;
        RECT 0.255 0.027 0.273 0.153 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.31 0.152 0.369 0.189 ;
        RECT 0.351 0.027 0.369 0.189 ;
        RECT 0.328 0.098 0.369 0.116 ;
        RECT 0.31 0.027 0.369 0.064 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.009 0.171 0.284 0.189 ;
        RECT 0.009 0.027 0.068 0.045 ;
        RECT 0.009 0.027 0.027 0.189 ;
    END
  END Y
END NAND5xp2R_ASAP7_6t_SL

MACRO NAND5xp2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND5xp2_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.063 0.119 0.081 ;
        RECT 0.045 0.135 0.113 0.153 ;
        RECT 0.045 0.063 0.063 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.144 0.027 0.162 0.146 ;
        RECT 0.088 0.099 0.162 0.117 ;
        RECT 0.099 0.027 0.162 0.045 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.027 0.23 0.068 ;
        RECT 0.18 0.135 0.227 0.153 ;
        RECT 0.18 0.027 0.198 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.252 0.115 0.291 0.153 ;
        RECT 0.252 0.027 0.289 0.066 ;
        RECT 0.234 0.098 0.27 0.116 ;
        RECT 0.252 0.027 0.27 0.153 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.309 0.151 0.36 0.189 ;
        RECT 0.342 0.027 0.36 0.189 ;
        RECT 0.319 0.098 0.36 0.116 ;
        RECT 0.31 0.027 0.36 0.066 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.009 0.171 0.284 0.189 ;
        RECT 0.009 0.027 0.068 0.045 ;
        RECT 0.009 0.027 0.027 0.189 ;
    END
  END Y
END NAND5xp2_ASAP7_6t_SL

MACRO NOR2x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.084 0.117 ;
        RECT 0.018 0.135 0.073 0.153 ;
        RECT 0.018 0.027 0.068 0.065 ;
        RECT 0.018 0.027 0.036 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.115 0.099 0.23 0.117 ;
        RECT 0.115 0.135 0.17 0.153 ;
        RECT 0.115 0.063 0.17 0.081 ;
        RECT 0.115 0.063 0.133 0.153 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.135 0.311 0.153 ;
        RECT 0.293 0.027 0.311 0.153 ;
        RECT 0.094 0.027 0.311 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.171 0.284 0.189 ;
  END
END NOR2x1_ASAP7_6t_SL

MACRO NOR2x2R_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2x2R_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.117 0.117 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.153 0.099 0.28 0.117 ;
        RECT 0.133 0.135 0.171 0.153 ;
        RECT 0.153 0.063 0.171 0.153 ;
        RECT 0.134 0.063 0.171 0.081 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.171 0.414 0.189 ;
        RECT 0.396 0.027 0.414 0.189 ;
        RECT 0.094 0.027 0.414 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.202 0.135 0.338 0.153 ;
      RECT 0.094 0.171 0.23 0.189 ;
  END
END NOR2x2R_ASAP7_6t_SL

MACRO NOR2x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.099 0.297 0.117 ;
        RECT 0.279 0.063 0.297 0.117 ;
        RECT 0.242 0.063 0.297 0.081 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.322 0.099 0.468 0.117 ;
        RECT 0.45 0.063 0.468 0.117 ;
        RECT 0.413 0.063 0.468 0.081 ;
        RECT 0.182 0.135 0.34 0.153 ;
        RECT 0.322 0.099 0.34 0.153 ;
        RECT 0.182 0.099 0.2 0.153 ;
        RECT 0.072 0.099 0.2 0.117 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.418 0.135 0.522 0.153 ;
        RECT 0.504 0.027 0.522 0.153 ;
        RECT 0.018 0.027 0.522 0.045 ;
        RECT 0.018 0.135 0.122 0.153 ;
        RECT 0.018 0.027 0.036 0.153 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.171 0.5 0.189 ;
  END
END NOR2x2_ASAP7_6t_SL

MACRO NOR2xp5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2xp5_ASAP7_6t_SL 0 0 ;
  SIZE 0.216 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.103 0.077 0.121 ;
        RECT 0.017 0.152 0.068 0.189 ;
        RECT 0.017 0.027 0.068 0.045 ;
        RECT 0.017 0.027 0.035 0.189 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.104 0.099 0.149 0.117 ;
        RECT 0.086 0.152 0.123 0.189 ;
        RECT 0.104 0.099 0.123 0.189 ;
        RECT 0.104 0.063 0.122 0.189 ;
        RECT 0.085 0.063 0.122 0.081 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.216 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.216 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.171 0.198 0.189 ;
        RECT 0.18 0.027 0.198 0.189 ;
        RECT 0.099 0.027 0.198 0.045 ;
    END
  END Y
END NOR2xp5_ASAP7_6t_SL

MACRO NOR3x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.594 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.099 0.468 0.117 ;
        RECT 0.45 0.063 0.468 0.117 ;
        RECT 0.396 0.063 0.468 0.081 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.133 0.099 0.338 0.117 ;
        RECT 0.133 0.135 0.225 0.153 ;
        RECT 0.133 0.027 0.177 0.071 ;
        RECT 0.133 0.027 0.151 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.079 0.117 ;
        RECT 0.018 0.027 0.073 0.045 ;
        RECT 0.018 0.147 0.068 0.189 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.594 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.418 0.171 0.576 0.189 ;
        RECT 0.558 0.027 0.576 0.189 ;
        RECT 0.202 0.027 0.576 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.256 0.135 0.5 0.153 ;
      RECT 0.094 0.171 0.338 0.189 ;
  END
END NOR3x1_ASAP7_6t_SL

MACRO NOR3x1f_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3x1f_ASAP7_6t_SL 0 0 ;
  SIZE 0.27 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.086 0.152 0.123 0.189 ;
        RECT 0.086 0.063 0.123 0.081 ;
        RECT 0.086 0.063 0.104 0.189 ;
        RECT 0.063 0.099 0.104 0.117 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.063 0.185 0.081 ;
        RECT 0.147 0.139 0.184 0.189 ;
        RECT 0.147 0.102 0.166 0.189 ;
        RECT 0.148 0.063 0.166 0.189 ;
        RECT 0.129 0.102 0.166 0.12 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.139 0.252 0.189 ;
        RECT 0.234 0.027 0.252 0.189 ;
        RECT 0.202 0.027 0.252 0.045 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.27 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.27 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.171 0.045 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END Y
END NOR3x1f_ASAP7_6t_SL

MACRO NOR3x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3x2_ASAP7_6t_SL 0 0 ;
  SIZE 1.08 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.946 0.099 1.001 0.117 ;
        RECT 0.983 0.063 1.001 0.117 ;
        RECT 0.153 0.063 1.001 0.081 ;
        RECT 0.094 0.099 0.171 0.117 ;
        RECT 0.153 0.063 0.171 0.117 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.519 0.135 0.579 0.153 ;
        RECT 0.519 0.099 0.575 0.117 ;
        RECT 0.519 0.099 0.537 0.153 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.08 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.08 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.88 0.171 1.062 0.189 ;
        RECT 1.044 0.027 1.062 0.189 ;
        RECT 0.018 0.027 1.062 0.045 ;
        RECT 0.018 0.171 0.176 0.189 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.31 0.099 0.752 0.117 ;
      LAYER M1 ;
        RECT 0.651 0.099 0.752 0.117 ;
        RECT 0.651 0.135 0.711 0.153 ;
        RECT 0.651 0.099 0.669 0.153 ;
        RECT 0.369 0.135 0.429 0.153 ;
        RECT 0.411 0.099 0.429 0.153 ;
        RECT 0.31 0.099 0.429 0.117 ;
      LAYER V1 ;
        RECT 0.315 0.099 0.333 0.117 ;
        RECT 0.729 0.099 0.747 0.117 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.742 0.135 0.986 0.153 ;
      RECT 0.256 0.171 0.824 0.189 ;
      RECT 0.094 0.135 0.338 0.153 ;
  END
END NOR3x2_ASAP7_6t_SL

MACRO NOR3xp33_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3xp33_ASAP7_6t_SL 0 0 ;
  SIZE 0.27 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.086 0.152 0.123 0.189 ;
        RECT 0.086 0.063 0.123 0.081 ;
        RECT 0.086 0.063 0.104 0.189 ;
        RECT 0.063 0.099 0.104 0.117 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.063 0.185 0.081 ;
        RECT 0.147 0.139 0.184 0.189 ;
        RECT 0.147 0.102 0.166 0.189 ;
        RECT 0.148 0.063 0.166 0.189 ;
        RECT 0.129 0.102 0.166 0.12 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.139 0.252 0.189 ;
        RECT 0.234 0.027 0.252 0.189 ;
        RECT 0.202 0.027 0.252 0.045 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.27 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.27 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.171 0.045 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END Y
END NOR3xp33_ASAP7_6t_SL

MACRO NOR4x3f_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4x3f_ASAP7_6t_SL 0 0 ;
  SIZE 0.756 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.575 0.099 0.645 0.117 ;
        RECT 0.627 0.063 0.645 0.117 ;
        RECT 0.487 0.063 0.645 0.081 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.353 0.099 0.501 0.117 ;
        RECT 0.353 0.063 0.396 0.153 ;
        RECT 0.264 0.063 0.396 0.081 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.153 0.099 0.29 0.117 ;
        RECT 0.093 0.135 0.171 0.153 ;
        RECT 0.153 0.063 0.171 0.153 ;
        RECT 0.094 0.063 0.171 0.081 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.117 0.117 ;
        RECT 0.018 0.027 0.068 0.065 ;
        RECT 0.018 0.149 0.067 0.189 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.756 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.756 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.171 0.738 0.189 ;
        RECT 0.72 0.027 0.738 0.189 ;
        RECT 0.094 0.027 0.738 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.092 0.171 0.216 0.189 ;
      RECT 0.198 0.135 0.216 0.189 ;
      RECT 0.198 0.135 0.328 0.153 ;
      RECT 0.428 0.135 0.666 0.153 ;
      RECT 0.25 0.171 0.5 0.189 ;
  END
END NOR4x3f_ASAP7_6t_SL

MACRO NOR4xp25_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4xp25_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.252 0.063 0.27 0.126 ;
        RECT 0.225 0.063 0.27 0.081 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.162 0.152 0.23 0.189 ;
        RECT 0.162 0.099 0.207 0.117 ;
        RECT 0.162 0.088 0.18 0.189 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.09 0.146 0.144 0.189 ;
        RECT 0.126 0.063 0.144 0.189 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.073 0.117 ;
        RECT 0.018 0.063 0.073 0.081 ;
        RECT 0.018 0.146 0.068 0.189 ;
        RECT 0.018 0.063 0.036 0.189 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.171 0.306 0.189 ;
        RECT 0.288 0.027 0.306 0.189 ;
        RECT 0.04 0.027 0.306 0.045 ;
    END
  END Y
END NOR4xp25_ASAP7_6t_SL

MACRO NOR5x1f_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR5x1f_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.171 0.074 0.189 ;
        RECT 0.018 0.043 0.036 0.189 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.105 0.171 0.144 0.189 ;
        RECT 0.126 0.063 0.144 0.189 ;
        RECT 0.098 0.063 0.144 0.081 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.162 0.15 0.217 0.189 ;
        RECT 0.162 0.063 0.217 0.102 ;
        RECT 0.18 0.063 0.198 0.189 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.235 0.063 0.312 0.081 ;
        RECT 0.235 0.171 0.293 0.189 ;
        RECT 0.235 0.063 0.253 0.189 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.324 0.171 0.361 0.189 ;
        RECT 0.343 0.027 0.361 0.189 ;
        RECT 0.324 0.027 0.361 0.045 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.055 0.027 0.285 0.045 ;
        RECT 0.055 0.135 0.096 0.153 ;
        RECT 0.055 0.027 0.073 0.153 ;
    END
  END Y
END NOR5x1f_ASAP7_6t_SL

MACRO NOR5xp2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR5xp2_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.135 0.119 0.153 ;
        RECT 0.045 0.063 0.113 0.081 ;
        RECT 0.045 0.063 0.063 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.171 0.162 0.189 ;
        RECT 0.144 0.07 0.162 0.189 ;
        RECT 0.088 0.099 0.162 0.117 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.148 0.23 0.189 ;
        RECT 0.18 0.063 0.227 0.081 ;
        RECT 0.18 0.063 0.198 0.189 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.252 0.063 0.291 0.101 ;
        RECT 0.252 0.15 0.289 0.189 ;
        RECT 0.252 0.063 0.27 0.189 ;
        RECT 0.234 0.1 0.27 0.118 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.31 0.15 0.36 0.189 ;
        RECT 0.342 0.027 0.36 0.189 ;
        RECT 0.319 0.1 0.36 0.118 ;
        RECT 0.309 0.027 0.36 0.065 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.009 0.027 0.284 0.045 ;
        RECT 0.009 0.171 0.068 0.189 ;
        RECT 0.009 0.027 0.027 0.189 ;
    END
  END Y
END NOR5xp2_ASAP7_6t_SL

MACRO O2A1O1A1Ixp33_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN O2A1O1A1Ixp33_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.171 0.055 0.189 ;
        RECT 0.018 0.063 0.055 0.081 ;
        RECT 0.018 0.063 0.036 0.189 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.105 0.099 0.144 0.117 ;
        RECT 0.086 0.135 0.123 0.153 ;
        RECT 0.105 0.064 0.123 0.153 ;
        RECT 0.086 0.064 0.123 0.082 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.135 0.218 0.153 ;
        RECT 0.18 0.063 0.218 0.081 ;
        RECT 0.18 0.063 0.198 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.287 0.135 0.325 0.153 ;
        RECT 0.287 0.063 0.325 0.081 ;
        RECT 0.287 0.063 0.305 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.135 0.414 0.153 ;
        RECT 0.396 0.064 0.414 0.153 ;
        RECT 0.376 0.064 0.414 0.082 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.171 0.468 0.189 ;
        RECT 0.45 0.027 0.468 0.189 ;
        RECT 0.423 0.027 0.468 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.207 0.027 0.387 0.045 ;
      RECT 0.099 0.171 0.225 0.189 ;
      RECT 0.04 0.027 0.171 0.045 ;
  END
END O2A1O1A1Ixp33_ASAP7_6t_SL

MACRO O2A1O1Ixp33_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN O2A1O1Ixp33_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.171 0.068 0.189 ;
        RECT 0.018 0.063 0.056 0.1 ;
        RECT 0.018 0.063 0.036 0.189 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1 0.099 0.142 0.117 ;
        RECT 0.081 0.135 0.118 0.153 ;
        RECT 0.1 0.063 0.118 0.153 ;
        RECT 0.081 0.063 0.118 0.1 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.154 0.135 0.195 0.153 ;
        RECT 0.177 0.063 0.195 0.153 ;
        RECT 0.154 0.063 0.195 0.081 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.249 0.063 0.267 0.136 ;
        RECT 0.215 0.116 0.252 0.153 ;
        RECT 0.22 0.063 0.267 0.081 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.171 0.315 0.189 ;
        RECT 0.297 0.027 0.315 0.189 ;
        RECT 0.207 0.027 0.315 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.099 0.171 0.225 0.189 ;
      RECT 0.04 0.027 0.171 0.045 ;
  END
END O2A1O1Ixp33_ASAP7_6t_SL

MACRO O2A1O1Ixp5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN O2A1O1Ixp5_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.232 0.063 0.25 0.104 ;
        RECT 0.018 0.063 0.25 0.081 ;
        RECT 0.018 0.027 0.117 0.045 ;
        RECT 0.018 0.171 0.068 0.189 ;
        RECT 0.018 0.027 0.037 0.081 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.085 0.099 0.176 0.117 ;
        RECT 0.085 0.099 0.122 0.153 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.296 0.063 0.344 0.081 ;
        RECT 0.291 0.064 0.309 0.122 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.331 0.135 0.38 0.153 ;
        RECT 0.362 0.094 0.38 0.153 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.398 0.027 0.416 0.157 ;
        RECT 0.315 0.027 0.416 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.256 0.171 0.333 0.189 ;
      RECT 0.256 0.135 0.274 0.189 ;
      RECT 0.153 0.135 0.274 0.153 ;
      RECT 0.148 0.027 0.284 0.045 ;
      RECT 0.099 0.171 0.225 0.189 ;
  END
END O2A1O1Ixp5_ASAP7_6t_SL

MACRO OA211x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA211x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.135 0.153 0.153 ;
        RECT 0.129 0.096 0.147 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.016 0.171 0.053 0.189 ;
        RECT 0.035 0.063 0.053 0.189 ;
        RECT 0.016 0.063 0.053 0.081 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.254 0.027 0.284 0.064 ;
        RECT 0.234 0.099 0.272 0.117 ;
        RECT 0.254 0.027 0.272 0.117 ;
        RECT 0.234 0.027 0.284 0.045 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.063 0.223 0.081 ;
        RECT 0.178 0.135 0.216 0.153 ;
        RECT 0.178 0.063 0.196 0.153 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.299 0.171 0.369 0.189 ;
        RECT 0.351 0.027 0.369 0.189 ;
        RECT 0.31 0.027 0.369 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.071 0.171 0.268 0.189 ;
      RECT 0.25 0.135 0.268 0.189 ;
      RECT 0.071 0.063 0.089 0.189 ;
      RECT 0.25 0.135 0.308 0.153 ;
      RECT 0.29 0.093 0.308 0.153 ;
      RECT 0.29 0.099 0.326 0.117 ;
      RECT 0.071 0.063 0.108 0.081 ;
      RECT 0.04 0.027 0.189 0.045 ;
  END
END OA211x1_ASAP7_6t_SL

MACRO OA211x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA211x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.135 0.153 0.153 ;
        RECT 0.129 0.09 0.147 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.016 0.171 0.053 0.189 ;
        RECT 0.035 0.063 0.053 0.189 ;
        RECT 0.016 0.063 0.053 0.081 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.254 0.027 0.31 0.076 ;
        RECT 0.234 0.099 0.272 0.117 ;
        RECT 0.254 0.027 0.272 0.117 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.135 0.265 0.153 ;
        RECT 0.178 0.063 0.223 0.081 ;
        RECT 0.178 0.063 0.196 0.153 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.328 0.171 0.412 0.189 ;
        RECT 0.394 0.027 0.412 0.189 ;
        RECT 0.328 0.027 0.412 0.045 ;
        RECT 0.328 0.147 0.346 0.189 ;
        RECT 0.328 0.027 0.346 0.068 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.071 0.171 0.309 0.189 ;
      RECT 0.291 0.099 0.309 0.189 ;
      RECT 0.071 0.063 0.089 0.189 ;
      RECT 0.291 0.099 0.346 0.117 ;
      RECT 0.071 0.063 0.108 0.081 ;
      RECT 0.035 0.027 0.193 0.045 ;
  END
END OA211x2_ASAP7_6t_SL

MACRO OA21x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.171 0.068 0.189 ;
        RECT 0.017 0.095 0.035 0.189 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.133 0.135 0.17 0.153 ;
        RECT 0.133 0.063 0.17 0.081 ;
        RECT 0.133 0.063 0.151 0.153 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.201 0.116 0.238 0.153 ;
        RECT 0.201 0.027 0.238 0.064 ;
        RECT 0.183 0.099 0.219 0.117 ;
        RECT 0.201 0.027 0.219 0.153 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.297 0.027 0.315 0.168 ;
        RECT 0.256 0.027 0.315 0.064 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.093 0.171 0.279 0.189 ;
      RECT 0.261 0.094 0.279 0.189 ;
      RECT 0.093 0.133 0.111 0.189 ;
      RECT 0.071 0.133 0.111 0.151 ;
      RECT 0.071 0.063 0.089 0.151 ;
      RECT 0.071 0.063 0.108 0.081 ;
      RECT 0.04 0.027 0.176 0.045 ;
  END
END OA21x1_ASAP7_6t_SL

MACRO OA21x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.016 0.171 0.068 0.189 ;
        RECT 0.016 0.095 0.034 0.189 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.133 0.135 0.17 0.153 ;
        RECT 0.133 0.063 0.17 0.081 ;
        RECT 0.133 0.063 0.151 0.153 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.201 0.116 0.238 0.153 ;
        RECT 0.201 0.027 0.238 0.045 ;
        RECT 0.182 0.099 0.219 0.117 ;
        RECT 0.201 0.027 0.219 0.153 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.293 0.027 0.351 0.045 ;
        RECT 0.263 0.135 0.311 0.153 ;
        RECT 0.293 0.027 0.311 0.153 ;
        RECT 0.258 0.063 0.311 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.093 0.171 0.359 0.189 ;
      RECT 0.341 0.094 0.359 0.189 ;
      RECT 0.093 0.133 0.111 0.189 ;
      RECT 0.071 0.133 0.111 0.151 ;
      RECT 0.071 0.063 0.09 0.151 ;
      RECT 0.071 0.063 0.108 0.081 ;
      RECT 0.04 0.027 0.171 0.045 ;
  END
END OA21x2_ASAP7_6t_SL

MACRO OA221x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA221x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.08 0.099 0.144 0.117 ;
        RECT 0.08 0.171 0.117 0.189 ;
        RECT 0.08 0.063 0.117 0.117 ;
        RECT 0.08 0.063 0.098 0.189 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.171 0.055 0.189 ;
        RECT 0.018 0.063 0.055 0.081 ;
        RECT 0.018 0.063 0.036 0.189 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.027 0.441 0.065 ;
        RECT 0.361 0.135 0.403 0.153 ;
        RECT 0.37 0.027 0.388 0.153 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.214 0.135 0.293 0.153 ;
        RECT 0.214 0.099 0.293 0.117 ;
        RECT 0.214 0.071 0.232 0.153 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.134 0.135 0.196 0.153 ;
        RECT 0.178 0.063 0.196 0.153 ;
        RECT 0.153 0.063 0.196 0.081 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.472 0.171 0.516 0.189 ;
        RECT 0.498 0.027 0.516 0.189 ;
        RECT 0.472 0.027 0.516 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.148 0.171 0.447 0.189 ;
      RECT 0.429 0.099 0.447 0.189 ;
      RECT 0.318 0.063 0.336 0.189 ;
      RECT 0.429 0.099 0.473 0.117 ;
      RECT 0.266 0.063 0.336 0.081 ;
      RECT 0.207 0.027 0.333 0.045 ;
      RECT 0.04 0.027 0.171 0.045 ;
  END
END OA221x1_ASAP7_6t_SL

MACRO OA221x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA221x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.594 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.08 0.099 0.144 0.117 ;
        RECT 0.08 0.171 0.117 0.189 ;
        RECT 0.08 0.063 0.117 0.117 ;
        RECT 0.08 0.063 0.098 0.189 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.171 0.055 0.189 ;
        RECT 0.018 0.063 0.055 0.081 ;
        RECT 0.018 0.063 0.036 0.189 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.027 0.441 0.065 ;
        RECT 0.361 0.135 0.403 0.153 ;
        RECT 0.37 0.027 0.388 0.153 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.214 0.135 0.293 0.153 ;
        RECT 0.214 0.099 0.293 0.117 ;
        RECT 0.214 0.071 0.232 0.153 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.134 0.135 0.196 0.153 ;
        RECT 0.178 0.063 0.196 0.153 ;
        RECT 0.153 0.063 0.196 0.081 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.594 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.472 0.171 0.551 0.189 ;
        RECT 0.531 0.027 0.551 0.189 ;
        RECT 0.472 0.027 0.551 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.148 0.171 0.447 0.189 ;
      RECT 0.429 0.099 0.447 0.189 ;
      RECT 0.318 0.063 0.336 0.189 ;
      RECT 0.429 0.099 0.473 0.117 ;
      RECT 0.266 0.063 0.336 0.081 ;
      RECT 0.207 0.027 0.333 0.045 ;
      RECT 0.04 0.027 0.171 0.045 ;
  END
END OA221x2_ASAP7_6t_SL

MACRO OA222x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA222x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.594 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.024 0.171 0.069 0.189 ;
        RECT 0.051 0.063 0.069 0.189 ;
        RECT 0.024 0.063 0.069 0.081 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.124 0.135 0.167 0.153 ;
        RECT 0.124 0.063 0.167 0.081 ;
        RECT 0.124 0.063 0.142 0.153 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.283 0.135 0.338 0.153 ;
        RECT 0.32 0.099 0.338 0.153 ;
        RECT 0.283 0.099 0.338 0.117 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.198 0.135 0.253 0.153 ;
        RECT 0.235 0.099 0.253 0.153 ;
        RECT 0.18 0.099 0.253 0.117 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.358 0.135 0.414 0.153 ;
        RECT 0.358 0.099 0.414 0.117 ;
        RECT 0.358 0.099 0.376 0.153 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.44 0.116 0.48 0.153 ;
        RECT 0.45 0.063 0.468 0.153 ;
        RECT 0.411 0.063 0.468 0.081 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.594 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.548 0.152 0.585 0.189 ;
        RECT 0.548 0.027 0.585 0.064 ;
        RECT 0.548 0.027 0.566 0.189 ;
        RECT 0.525 0.027 0.585 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.087 0.171 0.523 0.189 ;
      RECT 0.505 0.094 0.523 0.189 ;
      RECT 0.087 0.058 0.105 0.189 ;
      RECT 0.211 0.063 0.36 0.081 ;
      RECT 0.342 0.027 0.36 0.081 ;
      RECT 0.342 0.027 0.446 0.045 ;
      RECT 0.256 0.027 0.309 0.045 ;
      RECT 0.148 0.027 0.185 0.045 ;
      RECT 0.018 0.027 0.068 0.045 ;
    LAYER M2 ;
      RECT 0.04 0.027 0.287 0.045 ;
    LAYER V1 ;
      RECT 0.261 0.027 0.279 0.045 ;
      RECT 0.153 0.027 0.171 0.045 ;
      RECT 0.045 0.027 0.063 0.045 ;
  END
END OA222x1_ASAP7_6t_SL

MACRO OA222x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA222x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.648 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.016 0.099 0.07 0.117 ;
        RECT 0.052 0.076 0.07 0.117 ;
        RECT 0.016 0.152 0.068 0.189 ;
        RECT 0.016 0.099 0.034 0.189 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.124 0.135 0.167 0.153 ;
        RECT 0.124 0.063 0.162 0.081 ;
        RECT 0.124 0.063 0.142 0.153 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.283 0.135 0.338 0.153 ;
        RECT 0.32 0.099 0.338 0.153 ;
        RECT 0.283 0.099 0.338 0.117 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2 0.099 0.253 0.151 ;
        RECT 0.182 0.099 0.253 0.117 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.358 0.135 0.414 0.153 ;
        RECT 0.358 0.099 0.414 0.117 ;
        RECT 0.358 0.099 0.376 0.153 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.44 0.116 0.482 0.153 ;
        RECT 0.45 0.063 0.468 0.153 ;
        RECT 0.411 0.063 0.468 0.081 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.648 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.544 0.171 0.63 0.189 ;
        RECT 0.612 0.027 0.63 0.189 ;
        RECT 0.526 0.027 0.63 0.045 ;
        RECT 0.544 0.142 0.562 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.088 0.171 0.526 0.189 ;
      RECT 0.508 0.099 0.526 0.189 ;
      RECT 0.088 0.046 0.106 0.189 ;
      RECT 0.211 0.063 0.36 0.081 ;
      RECT 0.342 0.027 0.36 0.081 ;
      RECT 0.342 0.027 0.468 0.045 ;
      RECT 0.018 0.027 0.036 0.064 ;
      RECT 0.018 0.027 0.065 0.045 ;
      RECT 0.256 0.027 0.309 0.045 ;
      RECT 0.148 0.027 0.185 0.045 ;
    LAYER M2 ;
      RECT 0.02 0.027 0.287 0.045 ;
    LAYER V1 ;
      RECT 0.261 0.027 0.279 0.045 ;
      RECT 0.153 0.027 0.171 0.045 ;
      RECT 0.045 0.027 0.063 0.045 ;
  END
END OA222x2_ASAP7_6t_SL

MACRO OA22x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.031 0.171 0.068 0.189 ;
        RECT 0.05 0.063 0.068 0.189 ;
        RECT 0.031 0.063 0.068 0.081 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.105 0.1 0.141 0.118 ;
        RECT 0.086 0.152 0.123 0.189 ;
        RECT 0.105 0.063 0.123 0.189 ;
        RECT 0.086 0.063 0.123 0.1 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.309 0.135 0.346 0.153 ;
        RECT 0.309 0.027 0.346 0.045 ;
        RECT 0.309 0.027 0.327 0.153 ;
        RECT 0.291 0.099 0.327 0.117 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.151 0.192 0.189 ;
        RECT 0.174 0.063 0.192 0.189 ;
        RECT 0.155 0.063 0.192 0.081 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.418 0.171 0.458 0.189 ;
        RECT 0.44 0.027 0.458 0.189 ;
        RECT 0.418 0.027 0.458 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.235 0.171 0.393 0.189 ;
      RECT 0.375 0.099 0.393 0.189 ;
      RECT 0.235 0.063 0.254 0.189 ;
      RECT 0.217 0.144 0.254 0.162 ;
      RECT 0.375 0.099 0.415 0.117 ;
      RECT 0.217 0.063 0.254 0.081 ;
      RECT 0.04 0.027 0.284 0.045 ;
  END
END OA22x1_ASAP7_6t_SL

MACRO OA22x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.486 0.171 0.523 0.189 ;
        RECT 0.505 0.063 0.523 0.189 ;
        RECT 0.486 0.063 0.523 0.081 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.424 0.152 0.461 0.189 ;
        RECT 0.443 0.063 0.461 0.189 ;
        RECT 0.399 0.063 0.461 0.081 ;
        RECT 0.399 0.063 0.417 0.117 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.162 0.099 0.25 0.117 ;
        RECT 0.162 0.027 0.2 0.153 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.362 0.151 0.399 0.189 ;
        RECT 0.362 0.099 0.38 0.189 ;
        RECT 0.339 0.099 0.38 0.117 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.023 0.17 0.108 0.189 ;
        RECT 0.09 0.027 0.108 0.189 ;
        RECT 0.023 0.027 0.108 0.046 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.126 0.171 0.293 0.189 ;
      RECT 0.275 0.063 0.293 0.189 ;
      RECT 0.275 0.153 0.33 0.171 ;
      RECT 0.126 0.089 0.144 0.189 ;
      RECT 0.275 0.063 0.33 0.081 ;
      RECT 0.25 0.027 0.506 0.045 ;
  END
END OA22x2_ASAP7_6t_SL

MACRO OA311x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA311x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.135 0.217 0.153 ;
        RECT 0.18 0.094 0.198 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.144 0.189 ;
        RECT 0.126 0.063 0.144 0.189 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.101 0.093 0.119 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.063 0.252 0.122 ;
        RECT 0.215 0.063 0.252 0.081 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.269 0.135 0.306 0.153 ;
        RECT 0.288 0.07 0.306 0.153 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.472 0.171 0.521 0.189 ;
        RECT 0.503 0.027 0.521 0.189 ;
        RECT 0.472 0.027 0.521 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.198 0.171 0.36 0.189 ;
      RECT 0.342 0.027 0.36 0.189 ;
      RECT 0.342 0.099 0.473 0.117 ;
      RECT 0.31 0.027 0.36 0.045 ;
      RECT 0.094 0.027 0.234 0.045 ;
  END
END OA311x1_ASAP7_6t_SL

MACRO OA311x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA311x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.594 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.135 0.217 0.153 ;
        RECT 0.18 0.094 0.198 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.144 0.189 ;
        RECT 0.126 0.063 0.144 0.189 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.101 0.093 0.119 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.063 0.252 0.122 ;
        RECT 0.215 0.063 0.252 0.081 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.269 0.135 0.306 0.153 ;
        RECT 0.288 0.07 0.306 0.153 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.594 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.472 0.171 0.575 0.189 ;
        RECT 0.557 0.027 0.575 0.189 ;
        RECT 0.472 0.027 0.575 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.198 0.171 0.36 0.189 ;
      RECT 0.342 0.027 0.36 0.189 ;
      RECT 0.342 0.099 0.473 0.117 ;
      RECT 0.31 0.027 0.36 0.045 ;
      RECT 0.094 0.027 0.234 0.045 ;
  END
END OA311x2_ASAP7_6t_SL

MACRO OA31x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA31x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.115 0.116 0.153 0.153 ;
        RECT 0.123 0.063 0.141 0.153 ;
        RECT 0.098 0.063 0.141 0.081 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.135 0.222 0.153 ;
        RECT 0.174 0.063 0.211 0.081 ;
        RECT 0.178 0.063 0.196 0.153 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.255 0.027 0.292 0.064 ;
        RECT 0.231 0.099 0.273 0.117 ;
        RECT 0.255 0.027 0.273 0.117 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.171 0.054 0.189 ;
        RECT 0.017 0.058 0.035 0.189 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.305 0.171 0.36 0.189 ;
        RECT 0.342 0.027 0.36 0.189 ;
        RECT 0.323 0.027 0.36 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.079 0.171 0.274 0.189 ;
      RECT 0.256 0.135 0.274 0.189 ;
      RECT 0.079 0.124 0.097 0.189 ;
      RECT 0.256 0.135 0.324 0.153 ;
      RECT 0.306 0.094 0.324 0.153 ;
      RECT 0.055 0.124 0.097 0.142 ;
      RECT 0.055 0.058 0.073 0.142 ;
      RECT 0.094 0.027 0.23 0.045 ;
  END
END OA31x1_ASAP7_6t_SL

MACRO OA31x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA31x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.115 0.116 0.152 0.153 ;
        RECT 0.123 0.063 0.141 0.153 ;
        RECT 0.098 0.063 0.141 0.081 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.135 0.225 0.153 ;
        RECT 0.17 0.063 0.207 0.1 ;
        RECT 0.178 0.063 0.196 0.153 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.254 0.027 0.309 0.076 ;
        RECT 0.234 0.099 0.272 0.117 ;
        RECT 0.254 0.027 0.272 0.117 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.171 0.054 0.189 ;
        RECT 0.017 0.036 0.035 0.189 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.328 0.171 0.412 0.189 ;
        RECT 0.394 0.027 0.412 0.189 ;
        RECT 0.328 0.027 0.412 0.045 ;
        RECT 0.328 0.147 0.346 0.189 ;
        RECT 0.328 0.027 0.346 0.068 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.079 0.171 0.308 0.189 ;
      RECT 0.29 0.099 0.308 0.189 ;
      RECT 0.079 0.124 0.097 0.189 ;
      RECT 0.055 0.124 0.097 0.151 ;
      RECT 0.055 0.058 0.073 0.151 ;
      RECT 0.29 0.099 0.345 0.117 ;
      RECT 0.094 0.027 0.225 0.045 ;
  END
END OA31x2_ASAP7_6t_SL

MACRO OA321x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA321x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.594 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.594 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.094 0.198 0.146 ;
      LAYER M2 ;
        RECT 0.158 0.099 0.222 0.117 ;
      LAYER V1 ;
        RECT 0.18 0.099 0.198 0.117 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.144 0.189 ;
        RECT 0.126 0.063 0.144 0.189 ;
        RECT 0.098 0.063 0.144 0.081 ;
      LAYER M2 ;
        RECT 0.097 0.135 0.163 0.153 ;
      LAYER V1 ;
        RECT 0.126 0.135 0.144 0.153 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
      LAYER M2 ;
        RECT 0.018 0.099 0.082 0.117 ;
      LAYER V1 ;
        RECT 0.018 0.099 0.036 0.117 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.277 0.171 0.317 0.189 ;
        RECT 0.288 0.099 0.306 0.189 ;
      LAYER M2 ;
        RECT 0.257 0.135 0.336 0.153 ;
      LAYER V1 ;
        RECT 0.288 0.135 0.306 0.153 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.135 0.397 0.153 ;
        RECT 0.342 0.099 0.397 0.117 ;
        RECT 0.342 0.099 0.36 0.153 ;
      LAYER M2 ;
        RECT 0.328 0.099 0.403 0.117 ;
      LAYER V1 ;
        RECT 0.347 0.099 0.365 0.117 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.063 0.271 0.081 ;
        RECT 0.234 0.063 0.252 0.146 ;
      LAYER M2 ;
        RECT 0.212 0.063 0.278 0.081 ;
      LAYER V1 ;
        RECT 0.239 0.063 0.257 0.081 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.526 0.171 0.575 0.189 ;
        RECT 0.557 0.027 0.575 0.189 ;
        RECT 0.526 0.027 0.575 0.045 ;
      LAYER M2 ;
        RECT 0.372 0.027 0.575 0.045 ;
      LAYER V1 ;
        RECT 0.531 0.027 0.549 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.35 0.171 0.446 0.189 ;
      RECT 0.428 0.063 0.446 0.189 ;
      RECT 0.428 0.099 0.527 0.117 ;
      RECT 0.315 0.063 0.446 0.081 ;
      RECT 0.256 0.027 0.396 0.045 ;
      RECT 0.198 0.171 0.238 0.189 ;
      RECT 0.094 0.027 0.225 0.045 ;
    LAYER M2 ;
      RECT 0.207 0.171 0.441 0.189 ;
    LAYER V1 ;
      RECT 0.423 0.171 0.441 0.189 ;
      RECT 0.207 0.171 0.225 0.189 ;
  END
END OA321x1_ASAP7_6t_SL

MACRO OA321x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA321x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.648 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.648 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.094 0.198 0.146 ;
      LAYER M2 ;
        RECT 0.158 0.099 0.222 0.117 ;
      LAYER V1 ;
        RECT 0.18 0.099 0.198 0.117 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.144 0.189 ;
        RECT 0.126 0.063 0.144 0.189 ;
        RECT 0.107 0.063 0.144 0.081 ;
      LAYER M2 ;
        RECT 0.073 0.135 0.163 0.153 ;
      LAYER V1 ;
        RECT 0.126 0.135 0.144 0.153 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
      LAYER M2 ;
        RECT 0.018 0.099 0.082 0.117 ;
      LAYER V1 ;
        RECT 0.018 0.099 0.036 0.117 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.277 0.171 0.317 0.189 ;
        RECT 0.288 0.099 0.306 0.189 ;
      LAYER M2 ;
        RECT 0.257 0.135 0.336 0.153 ;
      LAYER V1 ;
        RECT 0.288 0.135 0.306 0.153 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.34 0.135 0.397 0.153 ;
        RECT 0.34 0.099 0.397 0.117 ;
        RECT 0.34 0.099 0.358 0.153 ;
      LAYER M2 ;
        RECT 0.33 0.099 0.403 0.117 ;
      LAYER V1 ;
        RECT 0.36 0.099 0.378 0.117 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.063 0.271 0.081 ;
        RECT 0.234 0.063 0.252 0.146 ;
      LAYER M2 ;
        RECT 0.212 0.063 0.278 0.081 ;
      LAYER V1 ;
        RECT 0.236 0.063 0.254 0.081 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.526 0.171 0.629 0.189 ;
        RECT 0.611 0.027 0.629 0.189 ;
        RECT 0.526 0.027 0.629 0.045 ;
      LAYER M2 ;
        RECT 0.459 0.099 0.629 0.117 ;
      LAYER V1 ;
        RECT 0.611 0.099 0.629 0.117 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.356 0.171 0.446 0.189 ;
      RECT 0.428 0.063 0.446 0.189 ;
      RECT 0.428 0.099 0.527 0.117 ;
      RECT 0.315 0.063 0.446 0.081 ;
      RECT 0.256 0.027 0.396 0.045 ;
      RECT 0.198 0.171 0.238 0.189 ;
      RECT 0.094 0.027 0.225 0.045 ;
    LAYER M2 ;
      RECT 0.207 0.171 0.441 0.189 ;
    LAYER V1 ;
      RECT 0.423 0.171 0.441 0.189 ;
      RECT 0.207 0.171 0.225 0.189 ;
  END
END OA321x2_ASAP7_6t_SL

MACRO OA322x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA322x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.648 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.537 0.063 0.559 0.137 ;
        RECT 0.518 0.152 0.555 0.189 ;
        RECT 0.537 0.063 0.555 0.189 ;
        RECT 0.504 0.099 0.559 0.117 ;
        RECT 0.522 0.063 0.559 0.117 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.152 0.5 0.189 ;
        RECT 0.45 0.063 0.487 0.081 ;
        RECT 0.45 0.063 0.468 0.189 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.359 0.063 0.425 0.081 ;
        RECT 0.364 0.171 0.414 0.189 ;
        RECT 0.396 0.063 0.414 0.189 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.208 0.135 0.267 0.153 ;
        RECT 0.249 0.099 0.267 0.153 ;
        RECT 0.209 0.099 0.267 0.117 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.285 0.099 0.361 0.117 ;
        RECT 0.285 0.135 0.34 0.153 ;
        RECT 0.285 0.099 0.303 0.153 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.152 0.068 0.189 ;
        RECT 0.017 0.063 0.054 0.189 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.122 0.099 0.178 0.117 ;
        RECT 0.122 0.135 0.177 0.153 ;
        RECT 0.122 0.099 0.14 0.153 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.648 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.171 0.631 0.189 ;
        RECT 0.613 0.037 0.631 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.577 0.027 0.595 0.122 ;
      RECT 0.526 0.027 0.595 0.045 ;
      RECT 0.086 0.171 0.333 0.189 ;
      RECT 0.086 0.101 0.104 0.189 ;
      RECT 0.072 0.027 0.091 0.119 ;
      RECT 0.032 0.027 0.091 0.045 ;
      RECT 0.109 0.063 0.328 0.081 ;
      RECT 0.109 0.04 0.127 0.081 ;
      RECT 0.261 0.027 0.495 0.045 ;
      RECT 0.193 0.027 0.23 0.045 ;
    LAYER M2 ;
      RECT 0.04 0.027 0.554 0.045 ;
    LAYER V1 ;
      RECT 0.531 0.027 0.549 0.045 ;
      RECT 0.207 0.027 0.225 0.045 ;
      RECT 0.045 0.027 0.063 0.045 ;
  END
END OA322x1_ASAP7_6t_SL

MACRO OA322x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA322x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.702 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.525 0.027 0.562 0.065 ;
        RECT 0.522 0.152 0.559 0.189 ;
        RECT 0.541 0.027 0.559 0.189 ;
        RECT 0.502 0.099 0.559 0.117 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.447 0.135 0.484 0.153 ;
        RECT 0.447 0.063 0.484 0.081 ;
        RECT 0.447 0.063 0.465 0.153 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.171 0.451 0.189 ;
        RECT 0.396 0.063 0.414 0.189 ;
        RECT 0.359 0.063 0.414 0.081 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.214 0.135 0.269 0.153 ;
        RECT 0.251 0.099 0.269 0.153 ;
        RECT 0.214 0.099 0.269 0.117 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.287 0.099 0.366 0.117 ;
        RECT 0.287 0.135 0.361 0.153 ;
        RECT 0.287 0.099 0.305 0.153 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.016 0.152 0.068 0.189 ;
        RECT 0.009 0.063 0.046 0.1 ;
        RECT 0.016 0.063 0.034 0.189 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.122 0.099 0.178 0.117 ;
        RECT 0.122 0.135 0.177 0.153 ;
        RECT 0.122 0.099 0.14 0.153 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.702 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.702 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.579 0.152 0.616 0.189 ;
        RECT 0.598 0.103 0.616 0.189 ;
        RECT 0.579 0.078 0.598 0.121 ;
        RECT 0.58 0.034 0.598 0.121 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.634 0.151 0.685 0.188 ;
      RECT 0.667 0.027 0.685 0.188 ;
      RECT 0.634 0.027 0.685 0.045 ;
      RECT 0.086 0.171 0.342 0.189 ;
      RECT 0.086 0.103 0.104 0.189 ;
      RECT 0.073 0.027 0.091 0.121 ;
      RECT 0.016 0.027 0.091 0.045 ;
      RECT 0.109 0.063 0.328 0.081 ;
      RECT 0.109 0.04 0.127 0.081 ;
      RECT 0.261 0.027 0.5 0.045 ;
      RECT 0.188 0.027 0.23 0.045 ;
    LAYER M2 ;
      RECT 0.035 0.027 0.683 0.045 ;
    LAYER V1 ;
      RECT 0.639 0.027 0.657 0.045 ;
      RECT 0.207 0.027 0.225 0.045 ;
      RECT 0.045 0.027 0.063 0.045 ;
  END
END OA322x2_ASAP7_6t_SL

MACRO OA32x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA32x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.214 0.137 0.251 0.174 ;
        RECT 0.233 0.063 0.251 0.174 ;
        RECT 0.214 0.063 0.251 0.1 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.159 0.137 0.196 0.174 ;
        RECT 0.178 0.063 0.196 0.174 ;
        RECT 0.159 0.063 0.196 0.1 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.123 0.063 0.141 0.151 ;
        RECT 0.099 0.063 0.141 0.081 ;
        RECT 0.085 0.027 0.122 0.064 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.09 0.306 0.174 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.379 0.132 0.416 0.152 ;
        RECT 0.398 0.063 0.416 0.152 ;
        RECT 0.36 0.063 0.416 0.1 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.023 0.027 0.06 0.045 ;
        RECT 0.023 0.027 0.041 0.175 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.324 0.171 0.393 0.189 ;
      RECT 0.324 0.056 0.342 0.189 ;
      RECT 0.064 0.171 0.12 0.189 ;
      RECT 0.064 0.099 0.082 0.189 ;
      RECT 0.363 0.027 0.416 0.045 ;
      RECT 0.153 0.027 0.287 0.045 ;
    LAYER M2 ;
      RECT 0.252 0.027 0.395 0.045 ;
      RECT 0.094 0.171 0.394 0.189 ;
    LAYER V1 ;
      RECT 0.369 0.027 0.387 0.045 ;
      RECT 0.369 0.171 0.387 0.189 ;
      RECT 0.261 0.027 0.279 0.045 ;
      RECT 0.099 0.171 0.117 0.189 ;
  END
END OA32x1_ASAP7_6t_SL

MACRO OA32x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA32x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.268 0.137 0.305 0.174 ;
        RECT 0.287 0.063 0.305 0.174 ;
        RECT 0.268 0.063 0.305 0.1 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.213 0.137 0.25 0.174 ;
        RECT 0.232 0.063 0.25 0.174 ;
        RECT 0.213 0.063 0.25 0.1 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.177 0.063 0.195 0.169 ;
        RECT 0.138 0.063 0.195 0.081 ;
        RECT 0.138 0.027 0.174 0.081 ;
        RECT 0.095 0.027 0.174 0.045 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.063 0.36 0.135 ;
        RECT 0.323 0.063 0.36 0.1 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.44 0.132 0.477 0.189 ;
        RECT 0.433 0.063 0.47 0.081 ;
        RECT 0.433 0.063 0.451 0.152 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.135 0.112 0.153 ;
        RECT 0.018 0.063 0.107 0.081 ;
        RECT 0.018 0.135 0.055 0.189 ;
        RECT 0.018 0.027 0.055 0.081 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.342 0.171 0.415 0.189 ;
      RECT 0.378 0.056 0.396 0.189 ;
      RECT 0.086 0.171 0.156 0.189 ;
      RECT 0.137 0.099 0.155 0.189 ;
      RECT 0.084 0.099 0.155 0.117 ;
      RECT 0.417 0.027 0.47 0.045 ;
      RECT 0.207 0.027 0.341 0.045 ;
    LAYER M2 ;
      RECT 0.31 0.027 0.446 0.045 ;
      RECT 0.091 0.171 0.392 0.189 ;
    LAYER V1 ;
      RECT 0.423 0.027 0.441 0.045 ;
      RECT 0.369 0.171 0.387 0.189 ;
      RECT 0.315 0.027 0.333 0.045 ;
      RECT 0.099 0.171 0.117 0.189 ;
  END
END OA32x2_ASAP7_6t_SL

MACRO OA331x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA331x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.063 0.271 0.081 ;
        RECT 0.224 0.171 0.261 0.189 ;
        RECT 0.234 0.063 0.252 0.189 ;
      LAYER M2 ;
        RECT 0.205 0.063 0.301 0.081 ;
      LAYER V1 ;
        RECT 0.247 0.063 0.265 0.081 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.171 0.063 0.208 0.081 ;
        RECT 0.162 0.171 0.199 0.189 ;
        RECT 0.181 0.063 0.199 0.189 ;
      LAYER M2 ;
        RECT 0.131 0.099 0.247 0.117 ;
      LAYER V1 ;
        RECT 0.181 0.099 0.199 0.117 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.063 0.144 0.12 ;
        RECT 0.107 0.063 0.144 0.081 ;
      LAYER M2 ;
        RECT 0.076 0.063 0.173 0.081 ;
      LAYER V1 ;
        RECT 0.117 0.063 0.135 0.081 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.286 0.171 0.323 0.189 ;
        RECT 0.286 0.099 0.304 0.189 ;
      LAYER M2 ;
        RECT 0.239 0.135 0.355 0.153 ;
      LAYER V1 ;
        RECT 0.286 0.135 0.304 0.153 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.334 0.099 0.371 0.117 ;
        RECT 0.343 0.099 0.361 0.146 ;
      LAYER M2 ;
        RECT 0.293 0.099 0.412 0.117 ;
      LAYER V1 ;
        RECT 0.347 0.099 0.365 0.117 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.135 0.443 0.153 ;
        RECT 0.396 0.106 0.414 0.153 ;
      LAYER M2 ;
        RECT 0.402 0.135 0.511 0.153 ;
      LAYER V1 ;
        RECT 0.423 0.135 0.441 0.153 ;
    END
  END B3
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.477 0.099 0.495 0.146 ;
        RECT 0.452 0.099 0.495 0.117 ;
      LAYER M2 ;
        RECT 0.446 0.099 0.511 0.117 ;
      LAYER V1 ;
        RECT 0.469 0.099 0.487 0.117 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.171 0.063 0.189 ;
        RECT 0.018 0.027 0.036 0.189 ;
      LAYER M2 ;
        RECT 0.039 0.027 0.137 0.045 ;
      LAYER V1 ;
        RECT 0.045 0.027 0.063 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.364 0.171 0.531 0.189 ;
      RECT 0.513 0.027 0.531 0.189 ;
      RECT 0.452 0.027 0.531 0.045 ;
      RECT 0.094 0.171 0.131 0.189 ;
      RECT 0.094 0.135 0.112 0.189 ;
      RECT 0.072 0.135 0.112 0.153 ;
      RECT 0.072 0.094 0.09 0.153 ;
      RECT 0.32 0.063 0.465 0.081 ;
      RECT 0.144 0.027 0.393 0.045 ;
    LAYER M2 ;
      RECT 0.094 0.171 0.446 0.189 ;
    LAYER V1 ;
      RECT 0.423 0.171 0.441 0.189 ;
      RECT 0.099 0.171 0.117 0.189 ;
  END
END OA331x1_ASAP7_6t_SL

MACRO OA331x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA331x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.594 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.594 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.063 0.327 0.081 ;
        RECT 0.288 0.063 0.306 0.163 ;
      LAYER M2 ;
        RECT 0.297 0.063 0.38 0.081 ;
      LAYER V1 ;
        RECT 0.297 0.063 0.315 0.081 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.225 0.063 0.262 0.081 ;
        RECT 0.233 0.063 0.251 0.163 ;
      LAYER M2 ;
        RECT 0.209 0.135 0.279 0.153 ;
      LAYER V1 ;
        RECT 0.233 0.135 0.251 0.153 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.063 0.198 0.119 ;
        RECT 0.161 0.063 0.198 0.081 ;
      LAYER M2 ;
        RECT 0.113 0.063 0.185 0.081 ;
      LAYER V1 ;
        RECT 0.167 0.063 0.185 0.081 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.336 0.099 0.364 0.117 ;
        RECT 0.34 0.099 0.358 0.163 ;
      LAYER M2 ;
        RECT 0.34 0.099 0.412 0.117 ;
      LAYER V1 ;
        RECT 0.34 0.099 0.358 0.117 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.383 0.135 0.425 0.153 ;
        RECT 0.397 0.106 0.415 0.153 ;
      LAYER M2 ;
        RECT 0.383 0.135 0.453 0.153 ;
      LAYER V1 ;
        RECT 0.388 0.135 0.406 0.153 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.135 0.534 0.153 ;
        RECT 0.45 0.106 0.468 0.153 ;
      LAYER M2 ;
        RECT 0.484 0.135 0.555 0.153 ;
      LAYER V1 ;
        RECT 0.484 0.135 0.502 0.153 ;
    END
  END B3
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.499 0.099 0.542 0.117 ;
      LAYER M2 ;
        RECT 0.5 0.099 0.572 0.117 ;
      LAYER V1 ;
        RECT 0.519 0.099 0.537 0.117 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.122 0.045 ;
        RECT 0.018 0.171 0.117 0.189 ;
        RECT 0.018 0.027 0.036 0.189 ;
      LAYER M2 ;
        RECT 0.018 0.027 0.256 0.045 ;
      LAYER V1 ;
        RECT 0.045 0.027 0.063 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.418 0.171 0.585 0.189 ;
      RECT 0.567 0.027 0.585 0.189 ;
      RECT 0.506 0.027 0.585 0.045 ;
      RECT 0.148 0.171 0.185 0.189 ;
      RECT 0.148 0.135 0.166 0.189 ;
      RECT 0.126 0.135 0.166 0.153 ;
      RECT 0.126 0.094 0.144 0.153 ;
      RECT 0.374 0.063 0.519 0.081 ;
      RECT 0.197 0.027 0.447 0.045 ;
    LAYER M2 ;
      RECT 0.153 0.171 0.466 0.189 ;
    LAYER V1 ;
      RECT 0.423 0.171 0.441 0.189 ;
      RECT 0.153 0.171 0.171 0.189 ;
  END
END OA331x2_ASAP7_6t_SL

MACRO OA332x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA332x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.756 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.159 0.101 0.2 0.119 ;
        RECT 0.094 0.171 0.177 0.189 ;
        RECT 0.159 0.058 0.177 0.189 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.068 0.135 0.141 0.153 ;
        RECT 0.123 0.063 0.141 0.153 ;
        RECT 0.094 0.063 0.141 0.081 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.171 0.055 0.189 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.171 0.249 0.189 ;
        RECT 0.231 0.063 0.249 0.189 ;
        RECT 0.212 0.063 0.249 0.081 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.267 0.171 0.338 0.189 ;
        RECT 0.267 0.099 0.322 0.117 ;
        RECT 0.267 0.099 0.285 0.189 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.31 0.135 0.412 0.153 ;
        RECT 0.357 0.099 0.412 0.117 ;
        RECT 0.357 0.099 0.375 0.153 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.592 0.135 0.632 0.153 ;
        RECT 0.614 0.027 0.632 0.153 ;
        RECT 0.58 0.027 0.632 0.045 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.445 0.135 0.53 0.153 ;
        RECT 0.512 0.099 0.53 0.153 ;
        RECT 0.445 0.099 0.53 0.117 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.756 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.756 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.701 0.171 0.738 0.189 ;
        RECT 0.72 0.027 0.738 0.189 ;
        RECT 0.688 0.027 0.738 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.369 0.171 0.668 0.189 ;
      RECT 0.65 0.099 0.668 0.189 ;
      RECT 0.549 0.063 0.567 0.189 ;
      RECT 0.65 0.099 0.695 0.117 ;
      RECT 0.482 0.063 0.567 0.081 ;
      RECT 0.275 0.063 0.451 0.081 ;
      RECT 0.433 0.027 0.451 0.081 ;
      RECT 0.433 0.027 0.549 0.045 ;
      RECT 0.193 0.027 0.392 0.045 ;
      RECT 0.094 0.027 0.135 0.045 ;
    LAYER M2 ;
      RECT 0.099 0.027 0.234 0.045 ;
    LAYER V1 ;
      RECT 0.207 0.027 0.225 0.045 ;
      RECT 0.099 0.027 0.117 0.045 ;
  END
END OA332x1_ASAP7_6t_SL

MACRO OA332x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA332x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.81 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.159 0.101 0.2 0.119 ;
        RECT 0.094 0.171 0.177 0.189 ;
        RECT 0.159 0.058 0.177 0.189 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.068 0.135 0.141 0.153 ;
        RECT 0.123 0.063 0.141 0.153 ;
        RECT 0.094 0.063 0.141 0.081 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.171 0.055 0.189 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.171 0.249 0.189 ;
        RECT 0.231 0.063 0.249 0.189 ;
        RECT 0.207 0.063 0.249 0.081 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.267 0.171 0.338 0.189 ;
        RECT 0.267 0.099 0.322 0.117 ;
        RECT 0.267 0.099 0.285 0.189 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.31 0.135 0.412 0.153 ;
        RECT 0.357 0.099 0.412 0.117 ;
        RECT 0.357 0.099 0.375 0.153 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.592 0.135 0.632 0.153 ;
        RECT 0.614 0.027 0.632 0.153 ;
        RECT 0.58 0.027 0.632 0.045 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.445 0.135 0.53 0.153 ;
        RECT 0.512 0.099 0.53 0.153 ;
        RECT 0.445 0.099 0.53 0.117 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.81 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.81 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.701 0.171 0.792 0.189 ;
        RECT 0.774 0.027 0.792 0.189 ;
        RECT 0.702 0.027 0.792 0.045 ;
        RECT 0.702 0.027 0.72 0.068 ;
        RECT 0.701 0.148 0.719 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.369 0.171 0.675 0.189 ;
      RECT 0.657 0.099 0.675 0.189 ;
      RECT 0.549 0.063 0.567 0.189 ;
      RECT 0.657 0.099 0.7 0.117 ;
      RECT 0.482 0.063 0.567 0.081 ;
      RECT 0.275 0.063 0.451 0.081 ;
      RECT 0.433 0.027 0.451 0.081 ;
      RECT 0.433 0.027 0.549 0.045 ;
      RECT 0.193 0.027 0.392 0.045 ;
      RECT 0.094 0.027 0.135 0.045 ;
    LAYER M2 ;
      RECT 0.099 0.027 0.234 0.045 ;
    LAYER V1 ;
      RECT 0.207 0.027 0.225 0.045 ;
      RECT 0.099 0.027 0.117 0.045 ;
  END
END OA332x2_ASAP7_6t_SL

MACRO OA333x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA333x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.864 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.684 0.135 0.721 0.153 ;
        RECT 0.684 0.063 0.721 0.081 ;
        RECT 0.684 0.063 0.702 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.629 0.063 0.666 0.153 ;
        RECT 0.556 0.099 0.666 0.117 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.171 0.638 0.189 ;
        RECT 0.58 0.135 0.598 0.189 ;
        RECT 0.466 0.135 0.598 0.153 ;
        RECT 0.466 0.099 0.521 0.117 ;
        RECT 0.466 0.099 0.484 0.153 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.171 0.249 0.189 ;
        RECT 0.231 0.063 0.249 0.189 ;
        RECT 0.205 0.063 0.249 0.081 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.267 0.171 0.322 0.189 ;
        RECT 0.267 0.099 0.322 0.117 ;
        RECT 0.267 0.057 0.285 0.189 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.357 0.099 0.417 0.117 ;
        RECT 0.31 0.135 0.412 0.153 ;
        RECT 0.357 0.099 0.375 0.153 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.159 0.101 0.2 0.119 ;
        RECT 0.094 0.171 0.177 0.189 ;
        RECT 0.159 0.058 0.177 0.189 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.093 0.135 0.141 0.153 ;
        RECT 0.123 0.063 0.141 0.153 ;
        RECT 0.094 0.063 0.141 0.081 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.864 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.864 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.796 0.171 0.846 0.189 ;
        RECT 0.828 0.027 0.846 0.189 ;
        RECT 0.796 0.027 0.846 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.688 0.171 0.764 0.189 ;
      RECT 0.746 0.132 0.764 0.189 ;
      RECT 0.757 0.066 0.775 0.15 ;
      RECT 0.746 0.027 0.764 0.084 ;
      RECT 0.634 0.027 0.764 0.045 ;
      RECT 0.313 0.063 0.603 0.081 ;
      RECT 0.585 0.04 0.603 0.081 ;
      RECT 0.313 0.04 0.331 0.081 ;
      RECT 0.505 0.027 0.554 0.045 ;
      RECT 0.364 0.171 0.549 0.189 ;
      RECT 0.363 0.027 0.413 0.045 ;
      RECT 0.193 0.027 0.239 0.045 ;
      RECT 0.094 0.027 0.135 0.045 ;
    LAYER M2 ;
      RECT 0.521 0.027 0.68 0.045 ;
      RECT 0.099 0.027 0.405 0.045 ;
    LAYER V1 ;
      RECT 0.639 0.027 0.657 0.045 ;
      RECT 0.531 0.027 0.549 0.045 ;
      RECT 0.369 0.027 0.387 0.045 ;
      RECT 0.207 0.027 0.225 0.045 ;
      RECT 0.099 0.027 0.117 0.045 ;
  END
END OA333x1_ASAP7_6t_SL

MACRO OA333x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA333x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.918 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.684 0.135 0.721 0.153 ;
        RECT 0.684 0.063 0.721 0.081 ;
        RECT 0.684 0.063 0.702 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.629 0.063 0.666 0.153 ;
        RECT 0.555 0.099 0.666 0.117 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.171 0.638 0.189 ;
        RECT 0.58 0.135 0.598 0.189 ;
        RECT 0.466 0.135 0.598 0.153 ;
        RECT 0.466 0.099 0.522 0.117 ;
        RECT 0.466 0.099 0.484 0.153 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.171 0.249 0.189 ;
        RECT 0.231 0.063 0.249 0.189 ;
        RECT 0.205 0.063 0.249 0.081 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.267 0.171 0.322 0.189 ;
        RECT 0.267 0.099 0.322 0.117 ;
        RECT 0.267 0.057 0.285 0.189 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.31 0.135 0.412 0.153 ;
        RECT 0.357 0.099 0.412 0.117 ;
        RECT 0.357 0.099 0.375 0.153 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.159 0.101 0.2 0.119 ;
        RECT 0.094 0.171 0.177 0.189 ;
        RECT 0.159 0.058 0.177 0.189 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.091 0.135 0.141 0.153 ;
        RECT 0.123 0.063 0.141 0.153 ;
        RECT 0.094 0.063 0.141 0.081 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.171 0.063 0.189 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.918 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.918 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.796 0.171 0.846 0.189 ;
        RECT 0.828 0.027 0.846 0.189 ;
        RECT 0.796 0.027 0.846 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.688 0.171 0.77 0.189 ;
      RECT 0.752 0.132 0.77 0.189 ;
      RECT 0.757 0.064 0.775 0.15 ;
      RECT 0.752 0.027 0.77 0.082 ;
      RECT 0.634 0.027 0.77 0.045 ;
      RECT 0.313 0.063 0.603 0.081 ;
      RECT 0.585 0.04 0.603 0.081 ;
      RECT 0.313 0.04 0.331 0.081 ;
      RECT 0.505 0.027 0.554 0.045 ;
      RECT 0.364 0.171 0.549 0.189 ;
      RECT 0.363 0.027 0.413 0.045 ;
      RECT 0.193 0.027 0.239 0.045 ;
      RECT 0.094 0.027 0.135 0.045 ;
    LAYER M2 ;
      RECT 0.521 0.027 0.68 0.045 ;
      RECT 0.099 0.027 0.405 0.045 ;
    LAYER V1 ;
      RECT 0.639 0.027 0.657 0.045 ;
      RECT 0.531 0.027 0.549 0.045 ;
      RECT 0.369 0.027 0.387 0.045 ;
      RECT 0.207 0.027 0.225 0.045 ;
      RECT 0.099 0.027 0.117 0.045 ;
  END
END OA333x2_ASAP7_6t_SL

MACRO OA33x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA33x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.152 0.252 0.189 ;
        RECT 0.234 0.063 0.252 0.189 ;
        RECT 0.187 0.063 0.252 0.081 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.277 0.063 0.317 0.081 ;
        RECT 0.277 0.135 0.315 0.153 ;
        RECT 0.288 0.063 0.306 0.153 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.137 0.099 0.203 0.117 ;
        RECT 0.137 0.171 0.176 0.189 ;
        RECT 0.137 0.046 0.155 0.189 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.28 0.171 0.358 0.189 ;
        RECT 0.34 0.106 0.358 0.189 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.171 0.458 0.189 ;
        RECT 0.376 0.099 0.417 0.117 ;
        RECT 0.376 0.099 0.394 0.189 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.485 0.171 0.524 0.189 ;
        RECT 0.485 0.099 0.522 0.117 ;
        RECT 0.485 0.099 0.503 0.189 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.071 0.143 0.112 0.161 ;
        RECT 0.071 0.063 0.112 0.081 ;
        RECT 0.02 0.171 0.089 0.189 ;
        RECT 0.071 0.063 0.089 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.426 0.135 0.467 0.153 ;
      RECT 0.449 0.063 0.467 0.153 ;
      RECT 0.353 0.063 0.504 0.081 ;
      RECT 0.472 0.027 0.504 0.081 ;
      RECT 0.472 0.027 0.522 0.045 ;
      RECT 0.018 0.027 0.036 0.124 ;
      RECT 0.018 0.027 0.073 0.045 ;
      RECT 0.201 0.027 0.441 0.045 ;
    LAYER M2 ;
      RECT 0.025 0.027 0.513 0.045 ;
    LAYER V1 ;
      RECT 0.477 0.027 0.495 0.045 ;
      RECT 0.045 0.027 0.063 0.045 ;
  END
END OA33x1_ASAP7_6t_SL

MACRO OA33x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA33x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.152 0.252 0.189 ;
        RECT 0.234 0.063 0.252 0.189 ;
        RECT 0.187 0.063 0.252 0.081 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.277 0.063 0.317 0.081 ;
        RECT 0.277 0.135 0.315 0.153 ;
        RECT 0.288 0.063 0.306 0.153 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.137 0.099 0.198 0.117 ;
        RECT 0.137 0.152 0.176 0.189 ;
        RECT 0.137 0.053 0.155 0.189 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.28 0.171 0.358 0.189 ;
        RECT 0.34 0.106 0.358 0.189 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.171 0.4455 0.189 ;
        RECT 0.376 0.099 0.417 0.117 ;
        RECT 0.376 0.099 0.394 0.189 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.488 0.135 0.531 0.189 ;
        RECT 0.506 0.099 0.524 0.189 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.071 0.143 0.112 0.161 ;
        RECT 0.089 0.058 0.107 0.112 ;
        RECT 0.02 0.171 0.089 0.189 ;
        RECT 0.071 0.094 0.089 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.426 0.135 0.467 0.153 ;
      RECT 0.449 0.063 0.467 0.153 ;
      RECT 0.353 0.063 0.497 0.081 ;
      RECT 0.474 0.027 0.497 0.081 ;
      RECT 0.474 0.027 0.522 0.045 ;
      RECT 0.018 0.027 0.036 0.124 ;
      RECT 0.018 0.027 0.068 0.046 ;
      RECT 0.201 0.027 0.441 0.045 ;
    LAYER M2 ;
      RECT 0.025 0.027 0.513 0.045 ;
    LAYER V1 ;
      RECT 0.477 0.027 0.495 0.045 ;
      RECT 0.045 0.027 0.063 0.045 ;
  END
END OA33x2_ASAP7_6t_SL

MACRO OAI211xp33_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211xp33_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.097 0.144 0.146 ;
      LAYER M2 ;
        RECT 0.096 0.099 0.17 0.117 ;
      LAYER V1 ;
        RECT 0.126 0.099 0.144 0.117 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.016 0.171 0.054 0.189 ;
        RECT 0.036 0.063 0.054 0.189 ;
        RECT 0.016 0.063 0.054 0.081 ;
      LAYER M2 ;
        RECT 0.018 0.135 0.115 0.153 ;
      LAYER V1 ;
        RECT 0.036 0.135 0.054 0.153 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.135 0.23 0.153 ;
        RECT 0.18 0.063 0.198 0.153 ;
        RECT 0.157 0.063 0.198 0.081 ;
      LAYER M2 ;
        RECT 0.135 0.063 0.223 0.081 ;
      LAYER V1 ;
        RECT 0.163 0.063 0.181 0.081 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.076 0.279 0.142 ;
        RECT 0.234 0.076 0.279 0.094 ;
        RECT 0.234 0.027 0.252 0.094 ;
        RECT 0.207 0.027 0.252 0.045 ;
      LAYER M2 ;
        RECT 0.218 0.099 0.295 0.117 ;
      LAYER V1 ;
        RECT 0.261 0.099 0.279 0.117 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.171 0.315 0.189 ;
        RECT 0.297 0.027 0.315 0.189 ;
        RECT 0.278 0.027 0.315 0.045 ;
        RECT 0.072 0.063 0.113 0.081 ;
        RECT 0.072 0.063 0.09 0.189 ;
      LAYER M2 ;
        RECT 0.156 0.171 0.308 0.189 ;
      LAYER V1 ;
        RECT 0.261 0.171 0.279 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.027 0.176 0.045 ;
  END
END OAI211xp33_ASAP7_6t_SL

MACRO OAI211xp67b_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211xp67b_ASAP7_6t_SL 0 0 ;
  SIZE 0.648 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.648 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.159 0.099 0.238 0.117 ;
        RECT 0.159 0.171 0.234 0.189 ;
        RECT 0.159 0.063 0.234 0.081 ;
        RECT 0.159 0.063 0.177 0.189 ;
      LAYER M2 ;
        RECT 0.168 0.099 0.232 0.117 ;
      LAYER V1 ;
        RECT 0.202 0.099 0.22 0.117 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.123 0.117 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
      LAYER M2 ;
        RECT 0.018 0.063 0.111 0.081 ;
      LAYER V1 ;
        RECT 0.018 0.063 0.036 0.081 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.314 0.171 0.369 0.189 ;
        RECT 0.314 0.099 0.369 0.117 ;
        RECT 0.314 0.099 0.332 0.189 ;
      LAYER M2 ;
        RECT 0.29 0.135 0.354 0.153 ;
      LAYER V1 ;
        RECT 0.314 0.135 0.332 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.526 0.171 0.564 0.189 ;
        RECT 0.546 0.099 0.564 0.189 ;
        RECT 0.519 0.099 0.564 0.117 ;
      LAYER M2 ;
        RECT 0.519 0.135 0.584 0.153 ;
      LAYER V1 ;
        RECT 0.546 0.135 0.564 0.153 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.583 0.171 0.631 0.189 ;
        RECT 0.583 0.063 0.603 0.189 ;
        RECT 0.519 0.063 0.603 0.081 ;
        RECT 0.418 0.171 0.495 0.189 ;
        RECT 0.094 0.171 0.131 0.189 ;
      LAYER M2 ;
        RECT 0.099 0.171 0.62 0.189 ;
      LAYER V1 ;
        RECT 0.099 0.171 0.117 0.189 ;
        RECT 0.423 0.171 0.441 0.189 ;
        RECT 0.585 0.171 0.603 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.288 0.063 0.449 0.081 ;
      RECT 0.288 0.027 0.306 0.081 ;
      RECT 0.094 0.027 0.306 0.045 ;
      RECT 0.361 0.027 0.608 0.045 ;
  END
END OAI211xp67b_ASAP7_6t_SL

MACRO OAI21xp25_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21xp25_ASAP7_6t_SL 0 0 ;
  SIZE 0.27 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.086 0.1 0.149 0.118 ;
        RECT 0.086 0.063 0.144 0.081 ;
        RECT 0.086 0.152 0.123 0.189 ;
        RECT 0.086 0.063 0.104 0.189 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.063 0.055 0.081 ;
        RECT 0.018 0.063 0.036 0.189 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.135 0.217 0.153 ;
        RECT 0.18 0.063 0.217 0.081 ;
        RECT 0.18 0.063 0.198 0.153 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.27 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.27 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.171 0.261 0.189 ;
        RECT 0.243 0.027 0.261 0.189 ;
        RECT 0.202 0.027 0.261 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.027 0.171 0.045 ;
  END
END OAI21xp25_ASAP7_6t_SL

MACRO OAI21xp5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21xp5_ASAP7_6t_SL 0 0 ;
  SIZE 0.27 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.086 0.1 0.144 0.118 ;
        RECT 0.086 0.063 0.144 0.081 ;
        RECT 0.086 0.1 0.123 0.189 ;
        RECT 0.086 0.063 0.104 0.189 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.148 0.068 0.189 ;
        RECT 0.018 0.063 0.061 0.081 ;
        RECT 0.018 0.063 0.036 0.189 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.135 0.217 0.153 ;
        RECT 0.18 0.063 0.217 0.081 ;
        RECT 0.18 0.063 0.198 0.153 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.27 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.27 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.171 0.261 0.189 ;
        RECT 0.243 0.027 0.261 0.189 ;
        RECT 0.202 0.027 0.261 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.027 0.171 0.045 ;
  END
END OAI21xp5_ASAP7_6t_SL

MACRO OAI21xp5b_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21xp5b_ASAP7_6t_SL 0 0 ;
  SIZE 0.27 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.016 0.171 0.053 0.189 ;
        RECT 0.035 0.063 0.053 0.189 ;
        RECT 0.016 0.063 0.053 0.081 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.145 0.063 0.196 0.153 ;
        RECT 0.122 0.1 0.196 0.118 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.214 0.171 0.251 0.189 ;
        RECT 0.214 0.027 0.251 0.045 ;
        RECT 0.214 0.027 0.232 0.189 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.27 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.27 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.071 0.171 0.177 0.189 ;
        RECT 0.071 0.063 0.114 0.081 ;
        RECT 0.071 0.063 0.089 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.027 0.176 0.045 ;
  END
END OAI21xp5b_ASAP7_6t_SL

MACRO OAI221xp33_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221xp33_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.264 0.063 0.301 0.081 ;
        RECT 0.254 0.099 0.282 0.182 ;
        RECT 0.264 0.063 0.282 0.182 ;
        RECT 0.234 0.099 0.282 0.117 ;
      LAYER M2 ;
        RECT 0.221 0.063 0.328 0.081 ;
      LAYER V1 ;
        RECT 0.275 0.063 0.293 0.081 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.332 0.063 0.369 0.1 ;
        RECT 0.307 0.171 0.362 0.189 ;
        RECT 0.344 0.063 0.362 0.189 ;
        RECT 0.307 0.135 0.362 0.153 ;
      LAYER M2 ;
        RECT 0.236 0.171 0.34 0.189 ;
      LAYER V1 ;
        RECT 0.315 0.171 0.333 0.189 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.009 0.152 0.047 0.189 ;
        RECT 0.016 0.134 0.047 0.189 ;
        RECT 0.009 0.063 0.047 0.1 ;
        RECT 0.016 0.063 0.034 0.189 ;
      LAYER M2 ;
        RECT 0.017 0.135 0.128 0.153 ;
      LAYER V1 ;
        RECT 0.022 0.135 0.04 0.153 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.101 0.099 0.147 0.117 ;
        RECT 0.101 0.099 0.12 0.146 ;
      LAYER M2 ;
        RECT 0.045 0.099 0.152 0.117 ;
      LAYER V1 ;
        RECT 0.124 0.099 0.142 0.117 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.135 0.217 0.153 ;
        RECT 0.159 0.063 0.217 0.081 ;
        RECT 0.18 0.063 0.198 0.153 ;
      LAYER M2 ;
        RECT 0.169 0.135 0.273 0.153 ;
      LAYER V1 ;
        RECT 0.182 0.135 0.2 0.153 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.065 0.171 0.225 0.189 ;
        RECT 0.065 0.063 0.12 0.081 ;
        RECT 0.065 0.063 0.083 0.189 ;
      LAYER M2 ;
        RECT 0.057 0.171 0.201 0.189 ;
      LAYER V1 ;
        RECT 0.099 0.171 0.117 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.207 0.027 0.362 0.045 ;
      RECT 0.04 0.027 0.171 0.045 ;
  END
END OAI221xp33_ASAP7_6t_SL

MACRO OAI221xp33f_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221xp33f_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.171 0.293 0.189 ;
        RECT 0.275 0.063 0.293 0.189 ;
        RECT 0.234 0.099 0.293 0.117 ;
        RECT 0.238 0.063 0.293 0.081 ;
      LAYER M2 ;
        RECT 0.235 0.063 0.304 0.081 ;
      LAYER V1 ;
        RECT 0.254 0.063 0.272 0.081 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.323 0.17 0.36 0.188 ;
        RECT 0.342 0.063 0.36 0.188 ;
        RECT 0.323 0.063 0.36 0.081 ;
      LAYER M2 ;
        RECT 0.291 0.099 0.36 0.117 ;
      LAYER V1 ;
        RECT 0.342 0.099 0.36 0.117 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.016 0.134 0.053 0.189 ;
        RECT 0.016 0.07 0.034 0.189 ;
      LAYER M2 ;
        RECT 0.016 0.099 0.085 0.117 ;
      LAYER V1 ;
        RECT 0.016 0.099 0.034 0.117 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.135 0.151 0.153 ;
        RECT 0.126 0.106 0.144 0.153 ;
      LAYER M2 ;
        RECT 0.11 0.135 0.174 0.153 ;
      LAYER V1 ;
        RECT 0.121 0.135 0.139 0.153 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.134 0.218 0.153 ;
        RECT 0.18 0.063 0.198 0.153 ;
        RECT 0.16 0.063 0.198 0.081 ;
      LAYER M2 ;
        RECT 0.157 0.099 0.226 0.117 ;
      LAYER V1 ;
        RECT 0.18 0.099 0.198 0.117 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.071 0.171 0.225 0.189 ;
        RECT 0.071 0.063 0.117 0.081 ;
        RECT 0.071 0.063 0.089 0.189 ;
      LAYER M2 ;
        RECT 0.071 0.063 0.194 0.081 ;
      LAYER V1 ;
        RECT 0.089 0.063 0.107 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.207 0.027 0.333 0.045 ;
      RECT 0.04 0.027 0.171 0.045 ;
  END
END OAI221xp33f_ASAP7_6t_SL

MACRO OAI222xp33_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222xp33_ASAP7_6t_SL 0 0 ;
  SIZE 0.54 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.54 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.54 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.009 0.132 0.046 0.189 ;
        RECT 0.018 0.07 0.036 0.189 ;
      LAYER M2 ;
        RECT 0.018 0.099 0.088 0.117 ;
      LAYER V1 ;
        RECT 0.018 0.099 0.036 0.117 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.128 0.099 0.157 0.117 ;
        RECT 0.109 0.135 0.146 0.153 ;
        RECT 0.128 0.099 0.146 0.153 ;
      LAYER M2 ;
        RECT 0.103 0.135 0.187 0.153 ;
      LAYER V1 ;
        RECT 0.115 0.135 0.133 0.153 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3 0.135 0.355 0.153 ;
        RECT 0.337 0.099 0.355 0.153 ;
        RECT 0.284 0.099 0.355 0.117 ;
      LAYER M2 ;
        RECT 0.287 0.135 0.371 0.153 ;
      LAYER V1 ;
        RECT 0.313 0.135 0.331 0.153 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.182 0.135 0.237 0.153 ;
        RECT 0.182 0.099 0.237 0.117 ;
        RECT 0.182 0.099 0.2 0.153 ;
      LAYER M2 ;
        RECT 0.164 0.099 0.26 0.117 ;
      LAYER V1 ;
        RECT 0.2 0.099 0.218 0.117 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.414 0.152 0.451 0.189 ;
        RECT 0.433 0.063 0.451 0.189 ;
        RECT 0.391 0.099 0.451 0.117 ;
        RECT 0.396 0.063 0.451 0.081 ;
      LAYER M2 ;
        RECT 0.365 0.099 0.461 0.117 ;
      LAYER V1 ;
        RECT 0.421 0.099 0.439 0.117 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.469 0.152 0.524 0.189 ;
        RECT 0.506 0.027 0.524 0.189 ;
        RECT 0.471 0.027 0.524 0.064 ;
      LAYER M2 ;
        RECT 0.405 0.063 0.524 0.081 ;
      LAYER V1 ;
        RECT 0.506 0.063 0.524 0.081 ;
    END
  END C2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.171 0.338 0.189 ;
        RECT 0.064 0.063 0.117 0.081 ;
        RECT 0.064 0.063 0.082 0.189 ;
      LAYER M2 ;
        RECT 0.069 0.063 0.187 0.081 ;
      LAYER V1 ;
        RECT 0.081 0.063 0.099 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.199 0.063 0.36 0.081 ;
      RECT 0.342 0.027 0.36 0.081 ;
      RECT 0.342 0.027 0.446 0.045 ;
      RECT 0.04 0.027 0.284 0.045 ;
  END
END OAI222xp33_ASAP7_6t_SL

MACRO OAI22xp5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22xp5_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.031 0.152 0.068 0.189 ;
        RECT 0.031 0.063 0.068 0.1 ;
        RECT 0.031 0.063 0.049 0.189 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.105 0.1 0.143 0.118 ;
        RECT 0.086 0.152 0.123 0.189 ;
        RECT 0.105 0.063 0.123 0.189 ;
        RECT 0.086 0.063 0.123 0.1 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.171 0.294 0.189 ;
        RECT 0.276 0.063 0.294 0.189 ;
        RECT 0.256 0.063 0.294 0.1 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.145 0.152 0.195 0.189 ;
        RECT 0.177 0.063 0.195 0.189 ;
        RECT 0.152 0.063 0.195 0.081 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.213 0.058 0.231 0.161 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.248 0.027 0.285 0.045 ;
      RECT 0.04 0.027 0.176 0.045 ;
    LAYER M2 ;
      RECT 0.148 0.027 0.284 0.045 ;
    LAYER V1 ;
      RECT 0.261 0.027 0.279 0.045 ;
      RECT 0.153 0.027 0.171 0.045 ;
  END
END OAI22xp5_ASAP7_6t_SL

MACRO OAI311xp33_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI311xp33_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.135 0.217 0.153 ;
        RECT 0.18 0.094 0.198 0.153 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.144 0.189 ;
        RECT 0.126 0.063 0.144 0.189 ;
        RECT 0.107 0.063 0.144 0.081 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.101 0.093 0.119 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.063 0.252 0.122 ;
        RECT 0.215 0.063 0.252 0.081 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.287 0.135 0.324 0.153 ;
        RECT 0.306 0.063 0.324 0.153 ;
        RECT 0.285 0.063 0.324 0.081 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.198 0.171 0.36 0.189 ;
        RECT 0.342 0.027 0.36 0.189 ;
        RECT 0.305 0.027 0.36 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.027 0.23 0.045 ;
  END
END OAI311xp33_ASAP7_6t_SL

MACRO OAI31x1f_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31x1f_ASAP7_6t_SL 0 0 ;
  SIZE 0.702 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.634 0.135 0.689 0.153 ;
        RECT 0.671 0.099 0.689 0.153 ;
        RECT 0.48 0.099 0.689 0.117 ;
        RECT 0.58 0.027 0.617 0.045 ;
        RECT 0.58 0.027 0.598 0.117 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.273 0.099 0.449 0.117 ;
        RECT 0.273 0.171 0.328 0.189 ;
        RECT 0.273 0.063 0.328 0.081 ;
        RECT 0.273 0.063 0.291 0.189 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.093 0.117 ;
        RECT 0.018 0.063 0.073 0.081 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.063 0.036 0.189 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.154 0.099 0.197 0.117 ;
        RECT 0.117 0.135 0.172 0.153 ;
        RECT 0.154 0.063 0.172 0.153 ;
        RECT 0.121 0.063 0.172 0.081 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.702 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.702 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.207 0.063 0.663 0.081 ;
      LAYER M1 ;
        RECT 0.629 0.063 0.674 0.081 ;
        RECT 0.201 0.171 0.255 0.189 ;
        RECT 0.237 0.063 0.255 0.189 ;
        RECT 0.207 0.063 0.255 0.081 ;
      LAYER V1 ;
        RECT 0.232 0.063 0.25 0.081 ;
        RECT 0.64 0.063 0.658 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.526 0.171 0.663 0.189 ;
      RECT 0.364 0.135 0.603 0.153 ;
      RECT 0.04 0.027 0.554 0.045 ;
      RECT 0.408 0.171 0.447 0.189 ;
      RECT 0.093 0.171 0.13 0.189 ;
    LAYER M2 ;
      RECT 0.094 0.171 0.447 0.189 ;
    LAYER V1 ;
      RECT 0.423 0.171 0.441 0.189 ;
      RECT 0.099 0.171 0.117 0.189 ;
  END
END OAI31x1f_ASAP7_6t_SL

MACRO OAI31xp5f_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31xp5f_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.154 0.135 0.195 0.153 ;
        RECT 0.177 0.063 0.195 0.153 ;
        RECT 0.154 0.063 0.195 0.081 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.105 0.1 0.141 0.118 ;
        RECT 0.086 0.152 0.123 0.189 ;
        RECT 0.105 0.063 0.123 0.189 ;
        RECT 0.086 0.063 0.123 0.081 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.062 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.22 0.135 0.257 0.153 ;
        RECT 0.239 0.063 0.257 0.153 ;
        RECT 0.22 0.063 0.257 0.081 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.183 0.171 0.306 0.189 ;
        RECT 0.288 0.056 0.306 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.093 0.027 0.239 0.045 ;
  END
END OAI31xp5f_ASAP7_6t_SL

MACRO OAI321xp33_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI321xp33_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.162 0.063 0.199 0.1 ;
        RECT 0.18 0.063 0.198 0.146 ;
      LAYER M2 ;
        RECT 0.158 0.099 0.222 0.117 ;
      LAYER V1 ;
        RECT 0.18 0.099 0.198 0.117 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.144 0.189 ;
        RECT 0.126 0.063 0.144 0.189 ;
        RECT 0.107 0.063 0.144 0.081 ;
      LAYER M2 ;
        RECT 0.097 0.135 0.163 0.153 ;
      LAYER V1 ;
        RECT 0.126 0.135 0.144 0.153 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.189 ;
      LAYER M2 ;
        RECT 0.018 0.063 0.105 0.081 ;
      LAYER V1 ;
        RECT 0.018 0.063 0.036 0.081 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.099 0.325 0.117 ;
        RECT 0.277 0.171 0.317 0.189 ;
        RECT 0.288 0.099 0.306 0.189 ;
      LAYER M2 ;
        RECT 0.268 0.099 0.347 0.117 ;
      LAYER V1 ;
        RECT 0.293 0.099 0.311 0.117 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.334 0.135 0.378 0.153 ;
        RECT 0.36 0.106 0.378 0.153 ;
      LAYER M2 ;
        RECT 0.336 0.135 0.403 0.153 ;
      LAYER V1 ;
        RECT 0.336 0.135 0.354 0.153 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.063 0.271 0.081 ;
        RECT 0.234 0.063 0.252 0.146 ;
      LAYER M2 ;
        RECT 0.212 0.063 0.278 0.081 ;
      LAYER V1 ;
        RECT 0.236 0.063 0.254 0.081 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.356 0.171 0.414 0.189 ;
        RECT 0.396 0.063 0.414 0.189 ;
        RECT 0.315 0.063 0.414 0.081 ;
        RECT 0.198 0.171 0.238 0.189 ;
      LAYER M2 ;
        RECT 0.207 0.171 0.387 0.189 ;
      LAYER V1 ;
        RECT 0.207 0.171 0.225 0.189 ;
        RECT 0.369 0.171 0.387 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.261 0.027 0.396 0.045 ;
      RECT 0.099 0.027 0.225 0.045 ;
  END
END OAI321xp33_ASAP7_6t_SL

MACRO OAI322xp33_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI322xp33_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.159 0.099 0.196 0.117 ;
        RECT 0.159 0.099 0.177 0.155 ;
      LAYER M2 ;
        RECT 0.141 0.099 0.22 0.117 ;
      LAYER V1 ;
        RECT 0.17 0.099 0.188 0.117 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.205 0.135 0.252 0.153 ;
        RECT 0.234 0.106 0.252 0.153 ;
      LAYER M2 ;
        RECT 0.202 0.135 0.27 0.153 ;
      LAYER V1 ;
        RECT 0.207 0.135 0.225 0.153 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.296 0.063 0.333 0.081 ;
        RECT 0.28 0.171 0.317 0.189 ;
        RECT 0.296 0.063 0.314 0.127 ;
        RECT 0.288 0.11 0.306 0.189 ;
      LAYER M2 ;
        RECT 0.271 0.063 0.362 0.081 ;
      LAYER V1 ;
        RECT 0.302 0.063 0.32 0.081 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.141 0.189 ;
        RECT 0.123 0.099 0.141 0.189 ;
        RECT 0.084 0.099 0.141 0.117 ;
      LAYER M2 ;
        RECT 0.076 0.135 0.153 0.153 ;
      LAYER V1 ;
        RECT 0.123 0.135 0.141 0.153 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.063 0.071 0.081 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.063 0.036 0.189 ;
      LAYER M2 ;
        RECT 0.018 0.063 0.097 0.081 ;
      LAYER V1 ;
        RECT 0.0365 0.063 0.0545 0.081 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.388 0.135 0.43 0.153 ;
        RECT 0.412 0.106 0.43 0.153 ;
      LAYER M2 ;
        RECT 0.378 0.135 0.448 0.153 ;
      LAYER V1 ;
        RECT 0.39 0.135 0.408 0.153 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.171 0.379 0.189 ;
        RECT 0.342 0.099 0.379 0.117 ;
        RECT 0.342 0.099 0.36 0.189 ;
      LAYER M2 ;
        RECT 0.326 0.099 0.4 0.117 ;
      LAYER V1 ;
        RECT 0.351 0.099 0.369 0.117 ;
    END
  END C2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.413 0.171 0.468 0.189 ;
        RECT 0.45 0.063 0.468 0.189 ;
        RECT 0.369 0.063 0.468 0.081 ;
        RECT 0.194 0.171 0.249 0.189 ;
      LAYER M2 ;
        RECT 0.202 0.171 0.446 0.189 ;
      LAYER V1 ;
        RECT 0.207 0.171 0.225 0.189 ;
        RECT 0.423 0.171 0.441 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.102 0.063 0.267 0.081 ;
      RECT 0.102 0.027 0.12 0.081 ;
      RECT 0.045 0.027 0.171 0.045 ;
      RECT 0.207 0.027 0.45 0.045 ;
  END
END OAI322xp33_ASAP7_6t_SL

MACRO OAI322xp33b_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI322xp33b_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.162 0.099 0.203 0.117 ;
        RECT 0.162 0.099 0.18 0.159 ;
      LAYER M2 ;
        RECT 0.15 0.099 0.214 0.117 ;
      LAYER V1 ;
        RECT 0.17 0.099 0.188 0.117 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.222 0.135 0.261 0.153 ;
        RECT 0.234 0.106 0.252 0.153 ;
      LAYER M2 ;
        RECT 0.207 0.135 0.283 0.153 ;
      LAYER V1 ;
        RECT 0.241 0.135 0.259 0.153 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.096 0.306 0.182 ;
      LAYER M2 ;
        RECT 0.247 0.099 0.311 0.117 ;
      LAYER V1 ;
        RECT 0.288 0.099 0.306 0.117 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.144 0.189 ;
        RECT 0.126 0.099 0.144 0.189 ;
        RECT 0.066 0.099 0.144 0.118 ;
      LAYER M2 ;
        RECT 0.089 0.135 0.171 0.153 ;
      LAYER V1 ;
        RECT 0.126 0.135 0.144 0.153 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.063 0.073 0.081 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.063 0.036 0.189 ;
      LAYER M2 ;
        RECT 0.018 0.063 0.09 0.081 ;
      LAYER V1 ;
        RECT 0.04 0.063 0.058 0.081 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.433 0.17 0.47 0.189 ;
        RECT 0.433 0.099 0.47 0.117 ;
        RECT 0.433 0.07 0.451 0.189 ;
      LAYER M2 ;
        RECT 0.404 0.135 0.468 0.153 ;
      LAYER V1 ;
        RECT 0.433 0.135 0.451 0.153 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.334 0.099 0.371 0.117 ;
        RECT 0.344 0.099 0.362 0.142 ;
      LAYER M2 ;
        RECT 0.342 0.099 0.406 0.117 ;
      LAYER V1 ;
        RECT 0.348 0.099 0.366 0.117 ;
    END
  END C2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.353 0.171 0.414 0.189 ;
        RECT 0.396 0.063 0.414 0.189 ;
        RECT 0.359 0.063 0.414 0.081 ;
        RECT 0.202 0.171 0.256 0.189 ;
      LAYER M2 ;
        RECT 0.207 0.171 0.387 0.189 ;
      LAYER V1 ;
        RECT 0.207 0.171 0.225 0.189 ;
        RECT 0.369 0.171 0.387 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.104 0.063 0.274 0.081 ;
      RECT 0.104 0.027 0.122 0.081 ;
      RECT 0.045 0.027 0.171 0.045 ;
      RECT 0.207 0.027 0.446 0.045 ;
  END
END OAI322xp33b_ASAP7_6t_SL

MACRO OAI32xp5f_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32xp5f_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.016 0.171 0.077 0.189 ;
        RECT 0.016 0.027 0.063 0.045 ;
        RECT 0.016 0.027 0.034 0.189 ;
      LAYER M2 ;
        RECT 0.038 0.171 0.168 0.189 ;
      LAYER V1 ;
        RECT 0.045 0.171 0.063 0.189 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.078 0.099 0.149 0.117 ;
      LAYER M2 ;
        RECT 0.061 0.099 0.163 0.117 ;
      LAYER V1 ;
        RECT 0.1 0.099 0.118 0.117 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.063 0.217 0.081 ;
        RECT 0.133 0.135 0.198 0.153 ;
        RECT 0.18 0.063 0.198 0.153 ;
      LAYER M2 ;
        RECT 0.147 0.063 0.249 0.081 ;
      LAYER V1 ;
        RECT 0.193 0.063 0.211 0.081 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.232 0.135 0.271 0.153 ;
        RECT 0.232 0.098 0.25 0.153 ;
      LAYER M2 ;
        RECT 0.215 0.135 0.307 0.153 ;
      LAYER V1 ;
        RECT 0.249 0.135 0.267 0.153 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.309 0.099 0.327 0.146 ;
        RECT 0.28 0.099 0.327 0.117 ;
      LAYER M2 ;
        RECT 0.243 0.099 0.345 0.117 ;
      LAYER V1 ;
        RECT 0.284 0.099 0.302 0.117 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.171 0.363 0.189 ;
        RECT 0.345 0.063 0.363 0.189 ;
        RECT 0.261 0.063 0.363 0.081 ;
        RECT 0.261 0.045 0.279 0.081 ;
      LAYER M2 ;
        RECT 0.209 0.171 0.338 0.189 ;
      LAYER V1 ;
        RECT 0.315 0.171 0.333 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.31 0.027 0.347 0.045 ;
      RECT 0.094 0.027 0.23 0.045 ;
    LAYER M2 ;
      RECT 0.148 0.027 0.338 0.045 ;
    LAYER V1 ;
      RECT 0.315 0.027 0.333 0.045 ;
      RECT 0.153 0.027 0.171 0.045 ;
  END
END OAI32xp5f_ASAP7_6t_SL

MACRO OAI331xp33_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI331xp33_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.063 0.224 0.081 ;
        RECT 0.18 0.063 0.198 0.146 ;
      LAYER M2 ;
        RECT 0.182 0.063 0.312 0.081 ;
      LAYER V1 ;
        RECT 0.2 0.063 0.218 0.081 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.155 0.189 ;
        RECT 0.094 0.063 0.155 0.081 ;
        RECT 0.126 0.063 0.144 0.189 ;
      LAYER M2 ;
        RECT 0.0865 0.135 0.1755 0.153 ;
      LAYER V1 ;
        RECT 0.126 0.135 0.144 0.153 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
      LAYER M2 ;
        RECT 0.039 0.027 0.128 0.045 ;
      LAYER V1 ;
        RECT 0.045 0.027 0.063 0.045 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.099 0.271 0.117 ;
        RECT 0.234 0.099 0.252 0.146 ;
      LAYER M2 ;
        RECT 0.153 0.099 0.311 0.117 ;
      LAYER V1 ;
        RECT 0.237 0.099 0.255 0.117 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.278 0.171 0.315 0.189 ;
        RECT 0.288 0.128 0.306 0.189 ;
      LAYER M2 ;
        RECT 0.207 0.135 0.311 0.153 ;
      LAYER V1 ;
        RECT 0.288 0.135 0.306 0.153 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.171 0.379 0.189 ;
        RECT 0.342 0.108 0.36 0.189 ;
      LAYER M2 ;
        RECT 0.342 0.135 0.42 0.153 ;
      LAYER V1 ;
        RECT 0.342 0.135 0.36 0.153 ;
    END
  END B3
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.412 0.076 0.43 0.146 ;
      LAYER M2 ;
        RECT 0.364 0.099 0.453 0.117 ;
      LAYER V1 ;
        RECT 0.412 0.099 0.43 0.117 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.41 0.171 0.468 0.189 ;
        RECT 0.45 0.027 0.468 0.189 ;
        RECT 0.418 0.027 0.468 0.045 ;
        RECT 0.195 0.171 0.237 0.189 ;
      LAYER M2 ;
        RECT 0.201 0.171 0.447 0.189 ;
      LAYER V1 ;
        RECT 0.207 0.171 0.225 0.189 ;
        RECT 0.423 0.171 0.441 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.261 0.063 0.387 0.081 ;
      RECT 0.369 0.035 0.387 0.081 ;
      RECT 0.099 0.027 0.333 0.045 ;
  END
END OAI331xp33_ASAP7_6t_SL

MACRO OAI332xp33_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI332xp33_ASAP7_6t_SL 0 0 ;
  SIZE 0.594 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.159 0.099 0.196 0.117 ;
        RECT 0.094 0.171 0.177 0.189 ;
        RECT 0.159 0.058 0.177 0.189 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.135 0.141 0.153 ;
        RECT 0.123 0.063 0.141 0.153 ;
        RECT 0.094 0.063 0.141 0.081 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.032 0.135 0.069 0.189 ;
        RECT 0.051 0.027 0.069 0.189 ;
        RECT 0.032 0.027 0.069 0.081 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.171 0.249 0.189 ;
        RECT 0.231 0.063 0.249 0.189 ;
        RECT 0.207 0.063 0.249 0.081 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.267 0.171 0.333 0.189 ;
        RECT 0.267 0.099 0.322 0.117 ;
        RECT 0.267 0.099 0.285 0.189 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.31 0.135 0.412 0.153 ;
        RECT 0.357 0.099 0.412 0.117 ;
        RECT 0.357 0.099 0.375 0.153 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.555 0.076 0.573 0.177 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.443 0.135 0.498 0.153 ;
        RECT 0.48 0.099 0.498 0.153 ;
        RECT 0.443 0.099 0.498 0.117 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.594 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.594 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.364 0.171 0.537 0.189 ;
        RECT 0.519 0.063 0.537 0.189 ;
        RECT 0.482 0.063 0.537 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.275 0.063 0.451 0.081 ;
      RECT 0.433 0.027 0.451 0.081 ;
      RECT 0.433 0.027 0.555 0.045 ;
      RECT 0.201 0.027 0.392 0.045 ;
      RECT 0.094 0.027 0.135 0.045 ;
    LAYER M2 ;
      RECT 0.094 0.027 0.234 0.045 ;
    LAYER V1 ;
      RECT 0.207 0.027 0.225 0.045 ;
      RECT 0.099 0.027 0.117 0.045 ;
  END
END OAI332xp33_ASAP7_6t_SL

MACRO OAI333xp33_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI333xp33_ASAP7_6t_SL 0 0 ;
  SIZE 0.702 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.171 0.656 0.189 ;
        RECT 0.638 0.087 0.656 0.189 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.559 0.135 0.617 0.153 ;
        RECT 0.599 0.099 0.617 0.153 ;
        RECT 0.559 0.099 0.617 0.117 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.448 0.099 0.522 0.117 ;
        RECT 0.448 0.135 0.521 0.153 ;
        RECT 0.448 0.099 0.466 0.153 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.171 0.255 0.189 ;
        RECT 0.237 0.1 0.255 0.189 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.291 0.135 0.346 0.153 ;
        RECT 0.328 0.099 0.346 0.153 ;
        RECT 0.291 0.099 0.346 0.117 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.375 0.135 0.43 0.153 ;
        RECT 0.412 0.099 0.43 0.153 ;
        RECT 0.375 0.099 0.43 0.117 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.063 0.23 0.081 ;
        RECT 0.159 0.128 0.196 0.149 ;
        RECT 0.178 0.063 0.196 0.149 ;
        RECT 0.094 0.171 0.177 0.189 ;
        RECT 0.159 0.128 0.177 0.189 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.104 0.135 0.141 0.153 ;
        RECT 0.123 0.063 0.141 0.153 ;
        RECT 0.094 0.063 0.141 0.081 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.032 0.135 0.069 0.189 ;
        RECT 0.051 0.027 0.069 0.189 ;
        RECT 0.032 0.027 0.069 0.081 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.702 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.702 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.521 0.027 0.68 0.045 ;
      LAYER M1 ;
        RECT 0.674 0.027 0.692 0.163 ;
        RECT 0.633 0.027 0.692 0.045 ;
        RECT 0.505 0.027 0.554 0.045 ;
      LAYER V1 ;
        RECT 0.531 0.027 0.549 0.045 ;
        RECT 0.639 0.027 0.657 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.265 0.063 0.603 0.081 ;
      RECT 0.585 0.04 0.603 0.081 ;
      RECT 0.265 0.04 0.283 0.081 ;
      RECT 0.315 0.171 0.549 0.189 ;
      RECT 0.315 0.027 0.393 0.045 ;
      RECT 0.094 0.027 0.23 0.045 ;
    LAYER M2 ;
      RECT 0.202 0.027 0.393 0.045 ;
    LAYER V1 ;
      RECT 0.369 0.027 0.387 0.045 ;
      RECT 0.207 0.027 0.225 0.045 ;
  END
END OAI333xp33_ASAP7_6t_SL

MACRO OAI33xp5f_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33xp5f_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.171 0.055 0.189 ;
        RECT 0.018 0.027 0.055 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.086 0.099 0.142 0.117 ;
        RECT 0.086 0.171 0.123 0.189 ;
        RECT 0.086 0.063 0.104 0.189 ;
        RECT 0.065 0.063 0.104 0.081 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.134 0.135 0.198 0.153 ;
        RECT 0.18 0.063 0.198 0.153 ;
        RECT 0.161 0.063 0.198 0.081 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.252 0.171 0.312 0.189 ;
        RECT 0.252 0.099 0.289 0.117 ;
        RECT 0.252 0.099 0.27 0.189 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.344 0.171 0.381 0.189 ;
        RECT 0.363 0.099 0.381 0.189 ;
        RECT 0.321 0.099 0.381 0.117 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.44 0.171 0.477 0.189 ;
        RECT 0.459 0.051 0.477 0.189 ;
        RECT 0.412 0.099 0.477 0.117 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.063 0.441 0.081 ;
        RECT 0.423 0.04 0.441 0.081 ;
        RECT 0.176 0.171 0.234 0.189 ;
        RECT 0.216 0.063 0.234 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.086 0.027 0.392 0.045 ;
  END
END OAI33xp5f_ASAP7_6t_SL

MACRO OR2x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.104 0.135 0.141 0.153 ;
        RECT 0.123 0.063 0.141 0.153 ;
        RECT 0.104 0.063 0.141 0.081 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.099 0.09 0.117 ;
        RECT 0.018 0.171 0.068 0.189 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.202 0.171 0.306 0.189 ;
        RECT 0.288 0.027 0.306 0.189 ;
        RECT 0.202 0.027 0.306 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.099 0.171 0.177 0.189 ;
      RECT 0.159 0.027 0.177 0.189 ;
      RECT 0.159 0.099 0.226 0.117 ;
      RECT 0.099 0.027 0.177 0.045 ;
  END
END OR2x2_ASAP7_6t_SL

MACRO OR2x3R_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2x3R_ASAP7_6t_SL 0 0 ;
  SIZE 0.648 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.153 0.063 0.171 0.11 ;
        RECT 0.018 0.063 0.171 0.081 ;
        RECT 0.018 0.171 0.069 0.189 ;
        RECT 0.018 0.063 0.036 0.189 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.215 0.099 0.257 0.117 ;
        RECT 0.094 0.135 0.234 0.153 ;
        RECT 0.215 0.099 0.234 0.153 ;
        RECT 0.094 0.135 0.131 0.189 ;
        RECT 0.094 0.099 0.112 0.189 ;
        RECT 0.072 0.099 0.112 0.117 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.648 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.648 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.315 0.171 0.63 0.189 ;
        RECT 0.612 0.027 0.63 0.189 ;
        RECT 0.287 0.027 0.63 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.202 0.171 0.284 0.189 ;
      RECT 0.266 0.135 0.284 0.189 ;
      RECT 0.266 0.135 0.306 0.153 ;
      RECT 0.288 0.063 0.306 0.153 ;
      RECT 0.234 0.063 0.306 0.081 ;
      RECT 0.234 0.027 0.252 0.081 ;
      RECT 0.094 0.027 0.252 0.045 ;
  END
END OR2x3R_ASAP7_6t_SL

MACRO OR2x4_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2x4_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.116 0.144 0.153 ;
        RECT 0.126 0.063 0.144 0.153 ;
        RECT 0.094 0.063 0.144 0.081 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.116 0.076 0.153 ;
        RECT 0.018 0.027 0.068 0.064 ;
        RECT 0.018 0.027 0.036 0.153 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.171 0.414 0.189 ;
        RECT 0.396 0.027 0.414 0.189 ;
        RECT 0.207 0.027 0.414 0.045 ;
        RECT 0.315 0.13 0.333 0.189 ;
        RECT 0.315 0.027 0.333 0.086 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.04 0.171 0.18 0.189 ;
      RECT 0.162 0.027 0.18 0.189 ;
      RECT 0.162 0.099 0.198 0.117 ;
      RECT 0.094 0.027 0.18 0.045 ;
  END
END OR2x4_ASAP7_6t_SL

MACRO OR3x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.324 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.063 0.055 0.081 ;
        RECT 0.018 0.063 0.036 0.189 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.107 0.099 0.144 0.117 ;
        RECT 0.088 0.152 0.125 0.189 ;
        RECT 0.107 0.063 0.125 0.189 ;
        RECT 0.088 0.063 0.125 0.081 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.161 0.135 0.198 0.153 ;
        RECT 0.18 0.063 0.198 0.153 ;
        RECT 0.161 0.063 0.198 0.081 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.324 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.324 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.171 0.306 0.189 ;
        RECT 0.288 0.027 0.306 0.189 ;
        RECT 0.261 0.027 0.306 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.153 0.171 0.234 0.189 ;
      RECT 0.216 0.027 0.234 0.189 ;
      RECT 0.216 0.099 0.262 0.117 ;
      RECT 0.04 0.027 0.234 0.045 ;
  END
END OR3x1_ASAP7_6t_SL

MACRO OR3x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.378 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.063 0.055 0.081 ;
        RECT 0.018 0.063 0.036 0.189 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.105 0.099 0.143 0.117 ;
        RECT 0.086 0.152 0.123 0.189 ;
        RECT 0.105 0.063 0.123 0.189 ;
        RECT 0.086 0.063 0.123 0.081 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.158 0.135 0.195 0.153 ;
        RECT 0.177 0.063 0.195 0.153 ;
        RECT 0.158 0.063 0.195 0.081 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.378 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.378 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.171 0.36 0.189 ;
        RECT 0.342 0.027 0.36 0.189 ;
        RECT 0.256 0.027 0.36 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.148 0.171 0.231 0.189 ;
      RECT 0.213 0.027 0.231 0.189 ;
      RECT 0.213 0.099 0.284 0.117 ;
      RECT 0.04 0.027 0.231 0.045 ;
  END
END OR3x2_ASAP7_6t_SL

MACRO OR3x4_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3x4_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.152 0.068 0.189 ;
        RECT 0.018 0.063 0.068 0.1 ;
        RECT 0.018 0.063 0.036 0.189 ;
      LAYER M2 ;
        RECT 0.018 0.063 0.089 0.081 ;
      LAYER V1 ;
        RECT 0.039 0.063 0.057 0.081 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.089 0.103 0.146 0.121 ;
        RECT 0.089 0.103 0.126 0.189 ;
      LAYER M2 ;
        RECT 0.067 0.135 0.172 0.153 ;
      LAYER V1 ;
        RECT 0.096 0.135 0.114 0.153 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.063 0.198 0.122 ;
        RECT 0.094 0.063 0.198 0.081 ;
      LAYER M2 ;
        RECT 0.15 0.099 0.224 0.117 ;
      LAYER V1 ;
        RECT 0.18 0.099 0.198 0.117 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.171 0.468 0.189 ;
        RECT 0.45 0.027 0.468 0.189 ;
        RECT 0.261 0.027 0.468 0.045 ;
        RECT 0.369 0.13 0.387 0.189 ;
        RECT 0.369 0.027 0.387 0.086 ;
      LAYER M2 ;
        RECT 0.348 0.099 0.468 0.117 ;
      LAYER V1 ;
        RECT 0.45 0.099 0.468 0.117 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.153 0.171 0.234 0.189 ;
      RECT 0.216 0.027 0.234 0.189 ;
      RECT 0.216 0.099 0.253 0.117 ;
      RECT 0.04 0.027 0.234 0.045 ;
  END
END OR3x4_ASAP7_6t_SL

MACRO OR4x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.009 0.151 0.063 0.188 ;
        RECT 0.009 0.027 0.063 0.064 ;
        RECT 0.009 0.099 0.047 0.117 ;
        RECT 0.009 0.027 0.027 0.188 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.081 0.099 0.144 0.117 ;
        RECT 0.081 0.152 0.118 0.189 ;
        RECT 0.081 0.063 0.118 0.117 ;
        RECT 0.081 0.063 0.099 0.189 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.136 0.135 0.198 0.153 ;
        RECT 0.18 0.063 0.198 0.153 ;
        RECT 0.16 0.063 0.198 0.081 ;
        RECT 0.136 0.135 0.173 0.189 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.227 0.135 0.264 0.153 ;
        RECT 0.227 0.063 0.264 0.081 ;
        RECT 0.235 0.063 0.253 0.153 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.325 0.171 0.392 0.189 ;
        RECT 0.325 0.027 0.392 0.045 ;
        RECT 0.325 0.027 0.343 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.207 0.171 0.307 0.189 ;
      RECT 0.289 0.027 0.307 0.189 ;
      RECT 0.094 0.027 0.307 0.045 ;
  END
END OR4x1_ASAP7_6t_SL

MACRO OR4x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.386 0.17 0.423 0.188 ;
        RECT 0.405 0.027 0.423 0.188 ;
        RECT 0.385 0.099 0.423 0.117 ;
        RECT 0.364 0.027 0.423 0.045 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.311 0.152 0.36 0.189 ;
        RECT 0.342 0.081 0.36 0.189 ;
        RECT 0.318 0.063 0.355 0.117 ;
        RECT 0.288 0.099 0.36 0.117 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.135 0.293 0.189 ;
        RECT 0.234 0.063 0.272 0.081 ;
        RECT 0.234 0.135 0.293 0.153 ;
        RECT 0.234 0.063 0.252 0.153 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.166 0.135 0.203 0.153 ;
        RECT 0.166 0.063 0.203 0.081 ;
        RECT 0.179 0.063 0.197 0.153 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.04 0.171 0.105 0.189 ;
        RECT 0.087 0.027 0.105 0.189 ;
        RECT 0.04 0.027 0.105 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.123 0.171 0.225 0.189 ;
      RECT 0.123 0.027 0.141 0.189 ;
      RECT 0.123 0.027 0.333 0.045 ;
  END
END OR4x2_ASAP7_6t_SL

MACRO OR5x1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR5x1_ASAP7_6t_SL 0 0 ;
  SIZE 0.432 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.016 0.171 0.065 0.189 ;
        RECT 0.016 0.043 0.034 0.189 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.097 0.171 0.141 0.189 ;
        RECT 0.123 0.063 0.141 0.189 ;
        RECT 0.103 0.063 0.141 0.081 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.171 0.227 0.189 ;
        RECT 0.178 0.063 0.196 0.189 ;
        RECT 0.159 0.063 0.196 0.1 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.252 0.164 0.289 0.189 ;
        RECT 0.252 0.132 0.27 0.189 ;
        RECT 0.231 0.132 0.27 0.15 ;
        RECT 0.214 0.063 0.251 0.1 ;
        RECT 0.231 0.063 0.249 0.15 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.321 0.126 0.339 0.182 ;
        RECT 0.295 0.063 0.334 0.081 ;
        RECT 0.295 0.126 0.339 0.144 ;
        RECT 0.295 0.063 0.313 0.144 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.432 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.432 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.367 0.171 0.416 0.189 ;
        RECT 0.398 0.052 0.416 0.189 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.071 0.107 0.089 0.15 ;
      RECT 0.052 0.107 0.089 0.125 ;
      RECT 0.359 0.027 0.377 0.114 ;
      RECT 0.052 0.027 0.07 0.125 ;
      RECT 0.052 0.027 0.377 0.045 ;
  END
END OR5x1_ASAP7_6t_SL

MACRO OR5x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR5x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.036 0.151 0.073 0.188 ;
        RECT 0.036 0.063 0.073 0.1 ;
        RECT 0.036 0.063 0.054 0.188 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.151 0.143 0.188 ;
        RECT 0.125 0.063 0.143 0.188 ;
        RECT 0.094 0.063 0.143 0.1 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.151 0.23 0.188 ;
        RECT 0.18 0.112 0.198 0.188 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.232 0.063 0.25 0.116 ;
        RECT 0.202 0.063 0.25 0.081 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.258 0.135 0.319 0.153 ;
        RECT 0.288 0.099 0.306 0.153 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.381 0.171 0.468 0.189 ;
        RECT 0.45 0.027 0.468 0.189 ;
        RECT 0.381 0.027 0.468 0.045 ;
        RECT 0.381 0.134 0.399 0.189 ;
        RECT 0.381 0.027 0.399 0.082 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.256 0.171 0.362 0.189 ;
      RECT 0.344 0.027 0.362 0.189 ;
      RECT 0.033 0.027 0.362 0.045 ;
  END
END OR5x2_ASAP7_6t_SL

MACRO SDFHx1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFHx1_ASAP7_6t_SL 0 0 ;
  SIZE 1.458 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.261 0.171 0.3 0.189 ;
        RECT 0.261 0.135 0.279 0.189 ;
        RECT 0.234 0.027 0.271 0.046 ;
        RECT 0.234 0.135 0.279 0.153 ;
        RECT 0.234 0.027 0.252 0.153 ;
      LAYER M2 ;
        RECT 0.135 0.135 0.358 0.153 ;
      LAYER V1 ;
        RECT 0.247 0.135 0.265 0.153 ;
    END
  END CLK
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.39 0.171 1.44 0.189 ;
        RECT 1.422 0.027 1.44 0.189 ;
        RECT 1.375 0.027 1.44 0.045 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.099 0.414 0.117 ;
        RECT 0.37 0.027 0.391 0.117 ;
        RECT 0.327 0.027 0.391 0.045 ;
        RECT 0.018 0.027 0.069 0.045 ;
        RECT 0.018 0.171 0.055 0.189 ;
        RECT 0.018 0.027 0.036 0.189 ;
      LAYER M2 ;
        RECT 0.02 0.027 0.398 0.045 ;
      LAYER V1 ;
        RECT 0.045 0.027 0.063 0.045 ;
        RECT 0.369 0.027 0.387 0.045 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.458 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.458 0.009 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.553 0.099 0.604 0.117 ;
      LAYER M2 ;
        RECT 0.502 0.099 0.632 0.117 ;
      LAYER V1 ;
        RECT 0.567 0.099 0.585 0.117 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.679 0.099 0.697 0.165 ;
        RECT 0.637 0.099 0.697 0.117 ;
      LAYER M2 ;
        RECT 0.663 0.099 0.793 0.117 ;
      LAYER V1 ;
        RECT 0.673 0.099 0.691 0.117 ;
    END
  END SI
  OBS
    LAYER M1 ;
      RECT 1.368 0.063 1.386 0.125 ;
      RECT 1.354 0.063 1.391 0.081 ;
      RECT 1.228 0.171 1.318 0.189 ;
      RECT 1.3 0.027 1.318 0.189 ;
      RECT 1.152 0.07 1.2 0.088 ;
      RECT 1.182 0.027 1.2 0.088 ;
      RECT 1.182 0.027 1.318 0.045 ;
      RECT 1.259 0.063 1.277 0.126 ;
      RECT 1.233 0.063 1.277 0.081 ;
      RECT 1.066 0.17 1.116 0.188 ;
      RECT 1.098 0.027 1.116 0.188 ;
      RECT 1.012 0.027 1.116 0.045 ;
      RECT 1.044 0.063 1.062 0.123 ;
      RECT 1.032 0.063 1.072 0.081 ;
      RECT 0.979 0.135 1.018 0.153 ;
      RECT 0.99 0.094 1.008 0.153 ;
      RECT 0.9 0.171 1.006 0.189 ;
      RECT 0.9 0.047 0.918 0.189 ;
      RECT 0.872 0.077 0.918 0.095 ;
      RECT 0.9 0.047 0.981 0.065 ;
      RECT 0.735 0.171 0.842 0.189 ;
      RECT 0.824 0.027 0.842 0.189 ;
      RECT 0.801 0.027 0.842 0.045 ;
      RECT 0.774 0.063 0.792 0.116 ;
      RECT 0.762 0.063 0.792 0.081 ;
      RECT 0.722 0.135 0.759 0.153 ;
      RECT 0.722 0.098 0.74 0.153 ;
      RECT 0.566 0.063 0.708 0.081 ;
      RECT 0.69 0.04 0.708 0.081 ;
      RECT 0.69 0.04 0.737 0.058 ;
      RECT 0.423 0.171 0.661 0.189 ;
      RECT 0.643 0.148 0.661 0.189 ;
      RECT 0.332 0.171 0.387 0.189 ;
      RECT 0.332 0.135 0.35 0.189 ;
      RECT 0.332 0.135 0.434 0.153 ;
      RECT 0.289 0.099 0.345 0.117 ;
      RECT 0.327 0.063 0.345 0.117 ;
      RECT 0.289 0.063 0.345 0.081 ;
      RECT 0.153 0.171 0.194 0.189 ;
      RECT 0.176 0.027 0.194 0.189 ;
      RECT 0.153 0.027 0.194 0.045 ;
      RECT 0.081 0.171 0.122 0.189 ;
      RECT 0.081 0.063 0.099 0.189 ;
      RECT 0.081 0.063 0.122 0.081 ;
      RECT 1.152 0.113 1.17 0.172 ;
      RECT 0.936 0.095 0.954 0.144 ;
      RECT 0.864 0.126 0.882 0.172 ;
      RECT 0.423 0.027 0.657 0.045 ;
      RECT 0.465 0.135 0.612 0.153 ;
      RECT 0.445 0.099 0.522 0.117 ;
    LAYER M2 ;
      RECT 1.098 0.063 1.391 0.081 ;
      RECT 0.396 0.135 1.17 0.153 ;
      RECT 0.153 0.063 1.062 0.081 ;
      RECT 0.824 0.099 0.954 0.117 ;
      RECT 0.073 0.099 0.47 0.117 ;
    LAYER V1 ;
      RECT 1.368 0.063 1.386 0.081 ;
      RECT 1.254 0.063 1.272 0.081 ;
      RECT 1.152 0.135 1.17 0.153 ;
      RECT 1.098 0.063 1.116 0.081 ;
      RECT 1.044 0.063 1.062 0.081 ;
      RECT 0.99 0.135 1.008 0.153 ;
      RECT 0.936 0.099 0.954 0.117 ;
      RECT 0.864 0.135 0.882 0.153 ;
      RECT 0.824 0.099 0.842 0.117 ;
      RECT 0.769 0.063 0.787 0.081 ;
      RECT 0.728 0.135 0.746 0.153 ;
      RECT 0.452 0.099 0.47 0.117 ;
      RECT 0.396 0.135 0.414 0.153 ;
      RECT 0.316 0.063 0.334 0.081 ;
      RECT 0.176 0.063 0.194 0.081 ;
      RECT 0.081 0.099 0.099 0.117 ;
  END
END SDFHx1_ASAP7_6t_SL

MACRO SDFHx2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFHx2_ASAP7_6t_SL 0 0 ;
  SIZE 1.512 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 1.206 0.171 1.326 0.189 ;
        RECT 1.308 0.027 1.326 0.189 ;
        RECT 1.282 0.027 1.326 0.046 ;
        RECT 1.206 0.094 1.224 0.189 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.33 0.099 0.385 0.117 ;
        RECT 0.33 0.062 0.348 0.117 ;
        RECT 0.287 0.062 0.348 0.081 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.39 0.171 1.44 0.189 ;
        RECT 1.422 0.027 1.44 0.189 ;
        RECT 1.375 0.027 1.44 0.045 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.099 0.185 0.117 ;
        RECT 0.032 0.171 0.166 0.189 ;
        RECT 0.148 0.099 0.166 0.189 ;
        RECT 0.032 0.027 0.069 0.045 ;
        RECT 0.032 0.027 0.05 0.189 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.418 0.171 0.484 0.189 ;
        RECT 0.466 0.099 0.484 0.189 ;
        RECT 0.418 0.099 0.484 0.117 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.512 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.512 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.242 0.135 1.283 0.153 ;
      RECT 1.242 0.051 1.26 0.153 ;
      RECT 1.152 0.051 1.17 0.122 ;
      RECT 1.152 0.051 1.26 0.069 ;
      RECT 0.972 0.171 1.04 0.189 ;
      RECT 0.972 0.027 0.99 0.189 ;
      RECT 0.935 0.07 0.99 0.088 ;
      RECT 0.972 0.027 1.04 0.045 ;
      RECT 0.85 0.17 0.91 0.188 ;
      RECT 0.892 0.027 0.91 0.188 ;
      RECT 0.796 0.027 0.91 0.045 ;
      RECT 0.828 0.063 0.846 0.123 ;
      RECT 0.816 0.063 0.856 0.081 ;
      RECT 0.763 0.135 0.802 0.153 ;
      RECT 0.774 0.094 0.792 0.153 ;
      RECT 0.684 0.171 0.79 0.189 ;
      RECT 0.684 0.047 0.702 0.189 ;
      RECT 0.666 0.077 0.702 0.095 ;
      RECT 0.684 0.047 0.765 0.065 ;
      RECT 0.531 0.171 0.626 0.189 ;
      RECT 0.608 0.027 0.626 0.189 ;
      RECT 0.585 0.027 0.626 0.045 ;
      RECT 0.556 0.063 0.574 0.116 ;
      RECT 0.537 0.063 0.574 0.081 ;
      RECT 0.366 0.063 0.501 0.081 ;
      RECT 0.483 0.027 0.501 0.081 ;
      RECT 0.366 0.04 0.384 0.081 ;
      RECT 0.483 0.027 0.549 0.045 ;
      RECT 0.507 0.135 0.544 0.153 ;
      RECT 0.507 0.102 0.525 0.153 ;
      RECT 0.207 0.135 0.225 0.178 ;
      RECT 0.207 0.135 0.441 0.153 ;
      RECT 0.086 0.135 0.123 0.153 ;
      RECT 0.086 0.063 0.105 0.153 ;
      RECT 0.228 0.099 0.299 0.117 ;
      RECT 0.228 0.063 0.246 0.117 ;
      RECT 0.086 0.063 0.246 0.081 ;
      RECT 1.368 0.088 1.386 0.125 ;
      RECT 1.116 0.058 1.134 0.158 ;
      RECT 1.008 0.089 1.026 0.126 ;
      RECT 0.935 0.113 0.953 0.172 ;
      RECT 0.72 0.095 0.738 0.144 ;
      RECT 0.648 0.126 0.666 0.172 ;
      RECT 0.415 0.027 0.452 0.045 ;
      RECT 0.261 0.171 0.387 0.189 ;
      RECT 0.198 0.027 0.235 0.045 ;
    LAYER M2 ;
      RECT 0.887 0.099 1.391 0.117 ;
      RECT 0.545 0.063 1.175 0.081 ;
      RECT 0.512 0.135 1.139 0.153 ;
      RECT 0.608 0.099 0.738 0.117 ;
      RECT 0.192 0.027 0.465 0.045 ;
    LAYER V1 ;
      RECT 1.368 0.099 1.386 0.117 ;
      RECT 1.152 0.063 1.17 0.081 ;
      RECT 1.116 0.135 1.134 0.153 ;
      RECT 1.008 0.099 1.026 0.117 ;
      RECT 0.935 0.135 0.953 0.153 ;
      RECT 0.892 0.099 0.91 0.117 ;
      RECT 0.828 0.063 0.846 0.081 ;
      RECT 0.774 0.135 0.792 0.153 ;
      RECT 0.72 0.099 0.738 0.117 ;
      RECT 0.648 0.135 0.666 0.153 ;
      RECT 0.608 0.099 0.626 0.117 ;
      RECT 0.55 0.063 0.568 0.081 ;
      RECT 0.517 0.135 0.535 0.153 ;
      RECT 0.423 0.027 0.441 0.045 ;
      RECT 0.207 0.027 0.225 0.045 ;
  END
END SDFHx2_ASAP7_6t_SL

MACRO SDFHx3_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFHx3_ASAP7_6t_SL 0 0 ;
  SIZE 1.566 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 1.206 0.171 1.326 0.189 ;
        RECT 1.308 0.027 1.326 0.189 ;
        RECT 1.282 0.027 1.326 0.046 ;
        RECT 1.206 0.094 1.224 0.189 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.33 0.099 0.385 0.117 ;
        RECT 0.33 0.062 0.348 0.117 ;
        RECT 0.287 0.062 0.348 0.081 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.39 0.171 1.548 0.189 ;
        RECT 1.53 0.027 1.548 0.189 ;
        RECT 1.375 0.027 1.548 0.045 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.099 0.185 0.117 ;
        RECT 0.032 0.171 0.166 0.189 ;
        RECT 0.148 0.099 0.166 0.189 ;
        RECT 0.032 0.027 0.069 0.045 ;
        RECT 0.032 0.027 0.05 0.189 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.418 0.171 0.484 0.189 ;
        RECT 0.466 0.099 0.484 0.189 ;
        RECT 0.418 0.099 0.484 0.117 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.566 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.566 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.242 0.135 1.283 0.153 ;
      RECT 1.242 0.051 1.26 0.153 ;
      RECT 1.152 0.051 1.17 0.122 ;
      RECT 1.152 0.051 1.26 0.069 ;
      RECT 0.972 0.171 1.04 0.189 ;
      RECT 0.972 0.027 0.99 0.189 ;
      RECT 0.935 0.07 0.99 0.088 ;
      RECT 0.972 0.027 1.04 0.045 ;
      RECT 0.85 0.17 0.91 0.188 ;
      RECT 0.892 0.027 0.91 0.188 ;
      RECT 0.796 0.027 0.91 0.045 ;
      RECT 0.828 0.063 0.846 0.123 ;
      RECT 0.816 0.063 0.856 0.081 ;
      RECT 0.763 0.135 0.802 0.153 ;
      RECT 0.774 0.094 0.792 0.153 ;
      RECT 0.684 0.171 0.79 0.189 ;
      RECT 0.684 0.047 0.702 0.189 ;
      RECT 0.666 0.077 0.702 0.095 ;
      RECT 0.684 0.047 0.765 0.065 ;
      RECT 0.531 0.171 0.626 0.189 ;
      RECT 0.608 0.027 0.626 0.189 ;
      RECT 0.585 0.027 0.626 0.045 ;
      RECT 0.556 0.063 0.574 0.116 ;
      RECT 0.537 0.063 0.574 0.081 ;
      RECT 0.366 0.063 0.501 0.081 ;
      RECT 0.483 0.027 0.501 0.081 ;
      RECT 0.366 0.04 0.384 0.081 ;
      RECT 0.483 0.027 0.549 0.045 ;
      RECT 0.507 0.135 0.544 0.153 ;
      RECT 0.507 0.102 0.525 0.153 ;
      RECT 0.207 0.135 0.225 0.178 ;
      RECT 0.207 0.135 0.441 0.153 ;
      RECT 0.086 0.135 0.123 0.153 ;
      RECT 0.086 0.063 0.105 0.153 ;
      RECT 0.228 0.099 0.299 0.117 ;
      RECT 0.228 0.063 0.246 0.117 ;
      RECT 0.086 0.063 0.246 0.081 ;
      RECT 1.358 0.099 1.502 0.117 ;
      RECT 1.116 0.058 1.134 0.158 ;
      RECT 1.008 0.089 1.026 0.126 ;
      RECT 0.935 0.113 0.953 0.172 ;
      RECT 0.72 0.095 0.738 0.144 ;
      RECT 0.648 0.126 0.666 0.172 ;
      RECT 0.415 0.027 0.452 0.045 ;
      RECT 0.261 0.171 0.387 0.189 ;
      RECT 0.198 0.027 0.235 0.045 ;
    LAYER M2 ;
      RECT 0.887 0.099 1.391 0.117 ;
      RECT 0.545 0.063 1.175 0.081 ;
      RECT 0.512 0.135 1.139 0.153 ;
      RECT 0.608 0.099 0.738 0.117 ;
      RECT 0.192 0.027 0.465 0.045 ;
    LAYER V1 ;
      RECT 1.368 0.099 1.386 0.117 ;
      RECT 1.152 0.063 1.17 0.081 ;
      RECT 1.116 0.135 1.134 0.153 ;
      RECT 1.008 0.099 1.026 0.117 ;
      RECT 0.935 0.135 0.953 0.153 ;
      RECT 0.892 0.099 0.91 0.117 ;
      RECT 0.828 0.063 0.846 0.081 ;
      RECT 0.774 0.135 0.792 0.153 ;
      RECT 0.72 0.099 0.738 0.117 ;
      RECT 0.648 0.135 0.666 0.153 ;
      RECT 0.608 0.099 0.626 0.117 ;
      RECT 0.55 0.063 0.568 0.081 ;
      RECT 0.517 0.135 0.535 0.153 ;
      RECT 0.423 0.027 0.441 0.045 ;
      RECT 0.207 0.027 0.225 0.045 ;
  END
END SDFHx3_ASAP7_6t_SL

MACRO SDFHx4_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFHx4_ASAP7_6t_SL 0 0 ;
  SIZE 1.62 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 1.206 0.171 1.326 0.189 ;
        RECT 1.308 0.027 1.326 0.189 ;
        RECT 1.282 0.027 1.326 0.046 ;
        RECT 1.206 0.094 1.224 0.189 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.33 0.099 0.385 0.117 ;
        RECT 0.33 0.062 0.348 0.117 ;
        RECT 0.287 0.062 0.348 0.081 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.39 0.171 1.576 0.189 ;
        RECT 1.558 0.027 1.576 0.189 ;
        RECT 1.39 0.027 1.576 0.045 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.099 0.185 0.117 ;
        RECT 0.032 0.171 0.166 0.189 ;
        RECT 0.148 0.099 0.166 0.189 ;
        RECT 0.032 0.027 0.069 0.045 ;
        RECT 0.032 0.027 0.05 0.189 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.418 0.171 0.484 0.189 ;
        RECT 0.466 0.099 0.484 0.189 ;
        RECT 0.418 0.099 0.484 0.117 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.62 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.62 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.242 0.135 1.283 0.153 ;
      RECT 1.242 0.051 1.26 0.153 ;
      RECT 1.152 0.051 1.17 0.122 ;
      RECT 1.152 0.051 1.26 0.069 ;
      RECT 0.972 0.171 1.04 0.189 ;
      RECT 0.972 0.027 0.99 0.189 ;
      RECT 0.935 0.07 0.99 0.088 ;
      RECT 0.972 0.027 1.04 0.045 ;
      RECT 0.85 0.17 0.91 0.188 ;
      RECT 0.892 0.027 0.91 0.188 ;
      RECT 0.796 0.027 0.91 0.045 ;
      RECT 0.828 0.063 0.846 0.123 ;
      RECT 0.816 0.063 0.856 0.081 ;
      RECT 0.763 0.135 0.802 0.153 ;
      RECT 0.774 0.094 0.792 0.153 ;
      RECT 0.684 0.171 0.79 0.189 ;
      RECT 0.684 0.047 0.702 0.189 ;
      RECT 0.666 0.077 0.702 0.095 ;
      RECT 0.684 0.047 0.765 0.065 ;
      RECT 0.531 0.171 0.626 0.189 ;
      RECT 0.608 0.027 0.626 0.189 ;
      RECT 0.585 0.027 0.626 0.045 ;
      RECT 0.556 0.063 0.574 0.116 ;
      RECT 0.537 0.063 0.574 0.081 ;
      RECT 0.366 0.063 0.501 0.081 ;
      RECT 0.483 0.027 0.501 0.081 ;
      RECT 0.366 0.04 0.384 0.081 ;
      RECT 0.483 0.027 0.549 0.045 ;
      RECT 0.507 0.135 0.544 0.153 ;
      RECT 0.507 0.102 0.525 0.153 ;
      RECT 0.207 0.135 0.225 0.178 ;
      RECT 0.207 0.135 0.441 0.153 ;
      RECT 0.086 0.135 0.123 0.153 ;
      RECT 0.086 0.063 0.105 0.153 ;
      RECT 0.228 0.099 0.299 0.117 ;
      RECT 0.228 0.063 0.246 0.117 ;
      RECT 0.086 0.063 0.246 0.081 ;
      RECT 1.363 0.099 1.526 0.117 ;
      RECT 1.116 0.058 1.134 0.158 ;
      RECT 1.008 0.089 1.026 0.126 ;
      RECT 0.935 0.113 0.953 0.172 ;
      RECT 0.72 0.095 0.738 0.144 ;
      RECT 0.648 0.126 0.666 0.172 ;
      RECT 0.415 0.027 0.452 0.045 ;
      RECT 0.261 0.171 0.387 0.189 ;
      RECT 0.198 0.027 0.235 0.045 ;
    LAYER M2 ;
      RECT 0.887 0.099 1.391 0.117 ;
      RECT 0.545 0.063 1.175 0.081 ;
      RECT 0.512 0.135 1.139 0.153 ;
      RECT 0.608 0.099 0.738 0.117 ;
      RECT 0.192 0.027 0.465 0.045 ;
    LAYER V1 ;
      RECT 1.368 0.099 1.386 0.117 ;
      RECT 1.152 0.063 1.17 0.081 ;
      RECT 1.116 0.135 1.134 0.153 ;
      RECT 1.008 0.099 1.026 0.117 ;
      RECT 0.935 0.135 0.953 0.153 ;
      RECT 0.892 0.099 0.91 0.117 ;
      RECT 0.828 0.063 0.846 0.081 ;
      RECT 0.774 0.135 0.792 0.153 ;
      RECT 0.72 0.099 0.738 0.117 ;
      RECT 0.648 0.135 0.666 0.153 ;
      RECT 0.608 0.099 0.626 0.117 ;
      RECT 0.55 0.063 0.568 0.081 ;
      RECT 0.517 0.135 0.535 0.153 ;
      RECT 0.423 0.027 0.441 0.045 ;
      RECT 0.207 0.027 0.225 0.045 ;
  END
END SDFHx4_ASAP7_6t_SL

MACRO SDFLx1_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFLx1_ASAP7_6t_SL 0 0 ;
  SIZE 1.458 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 1.206 0.171 1.326 0.189 ;
        RECT 1.308 0.027 1.326 0.189 ;
        RECT 1.282 0.027 1.326 0.046 ;
        RECT 1.206 0.094 1.224 0.189 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.33 0.099 0.385 0.117 ;
        RECT 0.33 0.062 0.348 0.117 ;
        RECT 0.287 0.062 0.348 0.081 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.39 0.171 1.44 0.189 ;
        RECT 1.422 0.027 1.44 0.189 ;
        RECT 1.385 0.027 1.44 0.045 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.099 0.185 0.117 ;
        RECT 0.032 0.171 0.166 0.189 ;
        RECT 0.148 0.099 0.166 0.189 ;
        RECT 0.032 0.027 0.069 0.045 ;
        RECT 0.032 0.027 0.05 0.189 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.418 0.171 0.484 0.189 ;
        RECT 0.466 0.099 0.484 0.189 ;
        RECT 0.418 0.099 0.484 0.117 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.458 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.458 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.152 0.051 1.17 0.158 ;
      RECT 1.242 0.135 1.283 0.153 ;
      RECT 1.242 0.051 1.26 0.153 ;
      RECT 1.152 0.051 1.26 0.069 ;
      RECT 0.972 0.171 1.04 0.189 ;
      RECT 0.972 0.027 0.99 0.189 ;
      RECT 0.935 0.07 0.99 0.088 ;
      RECT 0.972 0.027 1.04 0.045 ;
      RECT 0.85 0.17 0.91 0.188 ;
      RECT 0.892 0.027 0.91 0.188 ;
      RECT 0.796 0.027 0.91 0.045 ;
      RECT 0.828 0.063 0.846 0.123 ;
      RECT 0.816 0.063 0.856 0.081 ;
      RECT 0.763 0.135 0.802 0.153 ;
      RECT 0.774 0.094 0.792 0.153 ;
      RECT 0.684 0.171 0.79 0.189 ;
      RECT 0.684 0.047 0.702 0.189 ;
      RECT 0.666 0.077 0.702 0.095 ;
      RECT 0.684 0.047 0.765 0.065 ;
      RECT 0.531 0.171 0.626 0.189 ;
      RECT 0.608 0.027 0.626 0.189 ;
      RECT 0.585 0.027 0.626 0.045 ;
      RECT 0.556 0.063 0.574 0.116 ;
      RECT 0.537 0.063 0.574 0.081 ;
      RECT 0.366 0.063 0.501 0.081 ;
      RECT 0.483 0.027 0.501 0.081 ;
      RECT 0.366 0.04 0.384 0.081 ;
      RECT 0.483 0.027 0.549 0.045 ;
      RECT 0.507 0.135 0.544 0.153 ;
      RECT 0.507 0.102 0.525 0.153 ;
      RECT 0.207 0.135 0.225 0.178 ;
      RECT 0.207 0.135 0.441 0.153 ;
      RECT 0.086 0.135 0.123 0.153 ;
      RECT 0.086 0.063 0.105 0.153 ;
      RECT 0.228 0.099 0.299 0.117 ;
      RECT 0.228 0.063 0.246 0.117 ;
      RECT 0.086 0.063 0.246 0.081 ;
      RECT 1.368 0.088 1.386 0.125 ;
      RECT 1.116 0.058 1.134 0.158 ;
      RECT 1.008 0.089 1.026 0.126 ;
      RECT 0.935 0.113 0.953 0.172 ;
      RECT 0.72 0.095 0.738 0.144 ;
      RECT 0.648 0.126 0.666 0.172 ;
      RECT 0.415 0.027 0.452 0.045 ;
      RECT 0.261 0.171 0.387 0.189 ;
      RECT 0.198 0.027 0.235 0.045 ;
    LAYER M2 ;
      RECT 0.887 0.099 1.391 0.117 ;
      RECT 0.512 0.135 1.175 0.153 ;
      RECT 0.545 0.063 1.139 0.081 ;
      RECT 0.608 0.099 0.738 0.117 ;
      RECT 0.192 0.027 0.465 0.045 ;
    LAYER V1 ;
      RECT 1.368 0.099 1.386 0.117 ;
      RECT 1.152 0.135 1.17 0.153 ;
      RECT 1.116 0.063 1.134 0.081 ;
      RECT 1.008 0.099 1.026 0.117 ;
      RECT 0.935 0.135 0.953 0.153 ;
      RECT 0.892 0.099 0.91 0.117 ;
      RECT 0.828 0.063 0.846 0.081 ;
      RECT 0.774 0.135 0.792 0.153 ;
      RECT 0.72 0.099 0.738 0.117 ;
      RECT 0.648 0.135 0.666 0.153 ;
      RECT 0.608 0.099 0.626 0.117 ;
      RECT 0.55 0.063 0.568 0.081 ;
      RECT 0.517 0.135 0.535 0.153 ;
      RECT 0.423 0.027 0.441 0.045 ;
      RECT 0.207 0.027 0.225 0.045 ;
  END
END SDFLx1_ASAP7_6t_SL

MACRO SDFLx2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFLx2_ASAP7_6t_SL 0 0 ;
  SIZE 1.512 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 1.206 0.171 1.326 0.189 ;
        RECT 1.308 0.027 1.326 0.189 ;
        RECT 1.282 0.027 1.326 0.046 ;
        RECT 1.206 0.094 1.224 0.189 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.33 0.099 0.385 0.117 ;
        RECT 0.33 0.062 0.348 0.117 ;
        RECT 0.287 0.062 0.348 0.081 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.39 0.171 1.44 0.189 ;
        RECT 1.422 0.027 1.44 0.189 ;
        RECT 1.375 0.027 1.44 0.045 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.099 0.185 0.117 ;
        RECT 0.032 0.171 0.166 0.189 ;
        RECT 0.148 0.099 0.166 0.189 ;
        RECT 0.032 0.027 0.069 0.045 ;
        RECT 0.032 0.027 0.05 0.189 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.418 0.171 0.484 0.189 ;
        RECT 0.466 0.099 0.484 0.189 ;
        RECT 0.418 0.099 0.484 0.117 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.512 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.512 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.152 0.051 1.17 0.158 ;
      RECT 1.242 0.135 1.283 0.153 ;
      RECT 1.242 0.051 1.26 0.153 ;
      RECT 1.152 0.051 1.26 0.069 ;
      RECT 0.972 0.171 1.04 0.189 ;
      RECT 0.972 0.027 0.99 0.189 ;
      RECT 0.935 0.07 0.99 0.088 ;
      RECT 0.972 0.027 1.04 0.045 ;
      RECT 0.85 0.17 0.91 0.188 ;
      RECT 0.892 0.027 0.91 0.188 ;
      RECT 0.796 0.027 0.91 0.045 ;
      RECT 0.828 0.063 0.846 0.123 ;
      RECT 0.816 0.063 0.856 0.081 ;
      RECT 0.763 0.135 0.802 0.153 ;
      RECT 0.774 0.094 0.792 0.153 ;
      RECT 0.684 0.171 0.79 0.189 ;
      RECT 0.684 0.047 0.702 0.189 ;
      RECT 0.666 0.077 0.702 0.095 ;
      RECT 0.684 0.047 0.765 0.065 ;
      RECT 0.531 0.171 0.626 0.189 ;
      RECT 0.608 0.027 0.626 0.189 ;
      RECT 0.585 0.027 0.626 0.045 ;
      RECT 0.556 0.063 0.574 0.116 ;
      RECT 0.537 0.063 0.574 0.081 ;
      RECT 0.366 0.063 0.501 0.081 ;
      RECT 0.483 0.027 0.501 0.081 ;
      RECT 0.366 0.04 0.384 0.081 ;
      RECT 0.483 0.027 0.549 0.045 ;
      RECT 0.507 0.135 0.544 0.153 ;
      RECT 0.507 0.102 0.525 0.153 ;
      RECT 0.207 0.135 0.225 0.178 ;
      RECT 0.207 0.135 0.441 0.153 ;
      RECT 0.086 0.135 0.123 0.153 ;
      RECT 0.086 0.063 0.105 0.153 ;
      RECT 0.228 0.099 0.299 0.117 ;
      RECT 0.228 0.063 0.246 0.117 ;
      RECT 0.086 0.063 0.246 0.081 ;
      RECT 1.368 0.088 1.386 0.125 ;
      RECT 1.116 0.058 1.134 0.158 ;
      RECT 1.008 0.089 1.026 0.126 ;
      RECT 0.935 0.113 0.953 0.172 ;
      RECT 0.72 0.095 0.738 0.144 ;
      RECT 0.648 0.126 0.666 0.172 ;
      RECT 0.415 0.027 0.452 0.045 ;
      RECT 0.261 0.171 0.387 0.189 ;
      RECT 0.198 0.027 0.235 0.045 ;
    LAYER M2 ;
      RECT 0.887 0.099 1.391 0.117 ;
      RECT 0.512 0.135 1.175 0.153 ;
      RECT 0.545 0.063 1.139 0.081 ;
      RECT 0.608 0.099 0.738 0.117 ;
      RECT 0.192 0.027 0.465 0.045 ;
    LAYER V1 ;
      RECT 1.368 0.099 1.386 0.117 ;
      RECT 1.152 0.135 1.17 0.153 ;
      RECT 1.116 0.063 1.134 0.081 ;
      RECT 1.008 0.099 1.026 0.117 ;
      RECT 0.935 0.135 0.953 0.153 ;
      RECT 0.892 0.099 0.91 0.117 ;
      RECT 0.828 0.063 0.846 0.081 ;
      RECT 0.774 0.135 0.792 0.153 ;
      RECT 0.72 0.099 0.738 0.117 ;
      RECT 0.648 0.135 0.666 0.153 ;
      RECT 0.608 0.099 0.626 0.117 ;
      RECT 0.55 0.063 0.568 0.081 ;
      RECT 0.517 0.135 0.535 0.153 ;
      RECT 0.423 0.027 0.441 0.045 ;
      RECT 0.207 0.027 0.225 0.045 ;
  END
END SDFLx2_ASAP7_6t_SL

MACRO SDFLx3_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFLx3_ASAP7_6t_SL 0 0 ;
  SIZE 1.566 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 1.206 0.171 1.326 0.189 ;
        RECT 1.308 0.027 1.326 0.189 ;
        RECT 1.282 0.027 1.326 0.046 ;
        RECT 1.206 0.094 1.224 0.189 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.33 0.099 0.385 0.117 ;
        RECT 0.33 0.062 0.348 0.117 ;
        RECT 0.287 0.062 0.348 0.081 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.39 0.171 1.548 0.189 ;
        RECT 1.53 0.027 1.548 0.189 ;
        RECT 1.375 0.027 1.548 0.045 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.099 0.185 0.117 ;
        RECT 0.032 0.171 0.166 0.189 ;
        RECT 0.148 0.099 0.166 0.189 ;
        RECT 0.032 0.027 0.069 0.045 ;
        RECT 0.032 0.027 0.05 0.189 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.418 0.171 0.484 0.189 ;
        RECT 0.466 0.099 0.484 0.189 ;
        RECT 0.418 0.099 0.484 0.117 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.566 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.566 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.152 0.051 1.17 0.158 ;
      RECT 1.242 0.135 1.283 0.153 ;
      RECT 1.242 0.051 1.26 0.153 ;
      RECT 1.152 0.051 1.26 0.069 ;
      RECT 0.972 0.171 1.04 0.189 ;
      RECT 0.972 0.027 0.99 0.189 ;
      RECT 0.935 0.07 0.99 0.088 ;
      RECT 0.972 0.027 1.04 0.045 ;
      RECT 0.85 0.17 0.91 0.188 ;
      RECT 0.892 0.027 0.91 0.188 ;
      RECT 0.796 0.027 0.91 0.045 ;
      RECT 0.828 0.063 0.846 0.123 ;
      RECT 0.816 0.063 0.856 0.081 ;
      RECT 0.763 0.135 0.802 0.153 ;
      RECT 0.774 0.094 0.792 0.153 ;
      RECT 0.684 0.171 0.79 0.189 ;
      RECT 0.684 0.047 0.702 0.189 ;
      RECT 0.666 0.077 0.702 0.095 ;
      RECT 0.684 0.047 0.765 0.065 ;
      RECT 0.531 0.171 0.626 0.189 ;
      RECT 0.608 0.027 0.626 0.189 ;
      RECT 0.585 0.027 0.626 0.045 ;
      RECT 0.556 0.063 0.574 0.116 ;
      RECT 0.537 0.063 0.574 0.081 ;
      RECT 0.366 0.063 0.501 0.081 ;
      RECT 0.483 0.027 0.501 0.081 ;
      RECT 0.366 0.04 0.384 0.081 ;
      RECT 0.483 0.027 0.549 0.045 ;
      RECT 0.507 0.135 0.544 0.153 ;
      RECT 0.507 0.102 0.525 0.153 ;
      RECT 0.207 0.135 0.225 0.178 ;
      RECT 0.207 0.135 0.441 0.153 ;
      RECT 0.086 0.135 0.123 0.153 ;
      RECT 0.086 0.063 0.105 0.153 ;
      RECT 0.228 0.099 0.299 0.117 ;
      RECT 0.228 0.063 0.246 0.117 ;
      RECT 0.086 0.063 0.246 0.081 ;
      RECT 1.358 0.099 1.502 0.117 ;
      RECT 1.116 0.058 1.134 0.158 ;
      RECT 1.008 0.089 1.026 0.126 ;
      RECT 0.935 0.113 0.953 0.172 ;
      RECT 0.72 0.095 0.738 0.144 ;
      RECT 0.648 0.126 0.666 0.172 ;
      RECT 0.415 0.027 0.452 0.045 ;
      RECT 0.261 0.171 0.387 0.189 ;
      RECT 0.198 0.027 0.235 0.045 ;
    LAYER M2 ;
      RECT 0.887 0.099 1.391 0.117 ;
      RECT 0.512 0.135 1.175 0.153 ;
      RECT 0.545 0.063 1.139 0.081 ;
      RECT 0.608 0.099 0.738 0.117 ;
      RECT 0.192 0.027 0.465 0.045 ;
    LAYER V1 ;
      RECT 1.368 0.099 1.386 0.117 ;
      RECT 1.152 0.135 1.17 0.153 ;
      RECT 1.116 0.063 1.134 0.081 ;
      RECT 1.008 0.099 1.026 0.117 ;
      RECT 0.935 0.135 0.953 0.153 ;
      RECT 0.892 0.099 0.91 0.117 ;
      RECT 0.828 0.063 0.846 0.081 ;
      RECT 0.774 0.135 0.792 0.153 ;
      RECT 0.72 0.099 0.738 0.117 ;
      RECT 0.648 0.135 0.666 0.153 ;
      RECT 0.608 0.099 0.626 0.117 ;
      RECT 0.55 0.063 0.568 0.081 ;
      RECT 0.517 0.135 0.535 0.153 ;
      RECT 0.423 0.027 0.441 0.045 ;
      RECT 0.207 0.027 0.225 0.045 ;
  END
END SDFLx3_ASAP7_6t_SL

MACRO SDFLx4_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFLx4_ASAP7_6t_SL 0 0 ;
  SIZE 1.62 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 1.206 0.171 1.326 0.189 ;
        RECT 1.308 0.027 1.326 0.189 ;
        RECT 1.282 0.027 1.326 0.046 ;
        RECT 1.206 0.094 1.224 0.189 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.33 0.099 0.385 0.117 ;
        RECT 0.33 0.062 0.348 0.117 ;
        RECT 0.287 0.062 0.348 0.081 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.39 0.171 1.576 0.189 ;
        RECT 1.558 0.027 1.576 0.189 ;
        RECT 1.39 0.027 1.576 0.045 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.099 0.185 0.117 ;
        RECT 0.032 0.171 0.166 0.189 ;
        RECT 0.148 0.099 0.166 0.189 ;
        RECT 0.032 0.027 0.069 0.045 ;
        RECT 0.032 0.027 0.05 0.189 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.418 0.171 0.484 0.189 ;
        RECT 0.466 0.099 0.484 0.189 ;
        RECT 0.418 0.099 0.484 0.117 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 1.62 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.62 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.152 0.051 1.17 0.158 ;
      RECT 1.242 0.135 1.283 0.153 ;
      RECT 1.242 0.051 1.26 0.153 ;
      RECT 1.152 0.051 1.26 0.069 ;
      RECT 0.972 0.171 1.04 0.189 ;
      RECT 0.972 0.027 0.99 0.189 ;
      RECT 0.935 0.07 0.99 0.088 ;
      RECT 0.972 0.027 1.04 0.045 ;
      RECT 0.85 0.17 0.91 0.188 ;
      RECT 0.892 0.027 0.91 0.188 ;
      RECT 0.796 0.027 0.91 0.045 ;
      RECT 0.828 0.063 0.846 0.123 ;
      RECT 0.816 0.063 0.856 0.081 ;
      RECT 0.763 0.135 0.802 0.153 ;
      RECT 0.774 0.094 0.792 0.153 ;
      RECT 0.684 0.171 0.79 0.189 ;
      RECT 0.684 0.047 0.702 0.189 ;
      RECT 0.666 0.077 0.702 0.095 ;
      RECT 0.684 0.047 0.765 0.065 ;
      RECT 0.531 0.171 0.626 0.189 ;
      RECT 0.608 0.027 0.626 0.189 ;
      RECT 0.585 0.027 0.626 0.045 ;
      RECT 0.556 0.063 0.574 0.116 ;
      RECT 0.537 0.063 0.574 0.081 ;
      RECT 0.366 0.063 0.501 0.081 ;
      RECT 0.483 0.027 0.501 0.081 ;
      RECT 0.366 0.04 0.384 0.081 ;
      RECT 0.483 0.027 0.549 0.045 ;
      RECT 0.507 0.135 0.544 0.153 ;
      RECT 0.507 0.102 0.525 0.153 ;
      RECT 0.207 0.135 0.225 0.178 ;
      RECT 0.207 0.135 0.441 0.153 ;
      RECT 0.086 0.135 0.123 0.153 ;
      RECT 0.086 0.063 0.105 0.153 ;
      RECT 0.228 0.099 0.299 0.117 ;
      RECT 0.228 0.063 0.246 0.117 ;
      RECT 0.086 0.063 0.246 0.081 ;
      RECT 1.363 0.099 1.526 0.117 ;
      RECT 1.116 0.058 1.134 0.158 ;
      RECT 1.008 0.089 1.026 0.126 ;
      RECT 0.935 0.113 0.953 0.172 ;
      RECT 0.72 0.095 0.738 0.144 ;
      RECT 0.648 0.126 0.666 0.172 ;
      RECT 0.415 0.027 0.452 0.045 ;
      RECT 0.261 0.171 0.387 0.189 ;
      RECT 0.198 0.027 0.235 0.045 ;
    LAYER M2 ;
      RECT 0.887 0.099 1.391 0.117 ;
      RECT 0.512 0.135 1.175 0.153 ;
      RECT 0.545 0.063 1.139 0.081 ;
      RECT 0.608 0.099 0.738 0.117 ;
      RECT 0.192 0.027 0.465 0.045 ;
    LAYER V1 ;
      RECT 1.368 0.099 1.386 0.117 ;
      RECT 1.152 0.135 1.17 0.153 ;
      RECT 1.116 0.063 1.134 0.081 ;
      RECT 1.008 0.099 1.026 0.117 ;
      RECT 0.935 0.135 0.953 0.153 ;
      RECT 0.892 0.099 0.91 0.117 ;
      RECT 0.828 0.063 0.846 0.081 ;
      RECT 0.774 0.135 0.792 0.153 ;
      RECT 0.72 0.099 0.738 0.117 ;
      RECT 0.648 0.135 0.666 0.153 ;
      RECT 0.608 0.099 0.626 0.117 ;
      RECT 0.55 0.063 0.568 0.081 ;
      RECT 0.517 0.135 0.535 0.153 ;
      RECT 0.423 0.027 0.441 0.045 ;
      RECT 0.207 0.027 0.225 0.045 ;
  END
END SDFLx4_ASAP7_6t_SL

MACRO TAPCELL_ASAP7_6t_SL
  CLASS CORE WELLTAP ;
  ORIGIN 0 0 ;
  FOREIGN TAPCELL_ASAP7_6t_SL 0 0 ;
  SIZE 0.108 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.108 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.108 0.009 ;
    END
  END VSS
END TAPCELL_ASAP7_6t_SL

MACRO TAPCELL_WITH_FILLER_ASAP7_6t_SL
  CLASS CORE WELLTAP ;
  ORIGIN 0 0 ;
  FOREIGN TAPCELL_WITH_FILLER_ASAP7_6t_SL 0 0 ;
  SIZE 0.162 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.162 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.162 0.009 ;
    END
  END VSS
END TAPCELL_WITH_FILLER_ASAP7_6t_SL

MACRO TIEHIxp5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIEHIxp5_ASAP7_6t_SL 0 0 ;
  SIZE 0.162 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN H
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.144 0.189 ;
        RECT 0.126 0.027 0.144 0.189 ;
        RECT 0.067 0.072 0.144 0.09 ;
        RECT 0.094 0.027 0.144 0.045 ;
    END
  END H
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.162 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.162 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.018 0.128 0.095 0.146 ;
      RECT 0.018 0.027 0.036 0.146 ;
      RECT 0.018 0.027 0.063 0.045 ;
  END
END TIEHIxp5_ASAP7_6t_SL

MACRO TIELOxp5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIELOxp5_ASAP7_6t_SL 0 0 ;
  SIZE 0.162 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN L
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.171 0.144 0.189 ;
        RECT 0.126 0.027 0.144 0.189 ;
        RECT 0.067 0.126 0.144 0.144 ;
        RECT 0.094 0.027 0.144 0.045 ;
    END
  END L
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.162 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.162 0.009 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.018 0.171 0.063 0.189 ;
      RECT 0.018 0.07 0.036 0.189 ;
      RECT 0.018 0.07 0.095 0.088 ;
  END
END TIELOxp5_ASAP7_6t_SL

MACRO XNOR2x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.702 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.056 0.099 0.144 0.117 ;
        RECT 0.08 0.063 0.122 0.117 ;
        RECT 0.056 0.072 0.095 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.099 0.36 0.117 ;
        RECT 0.018 0.171 0.225 0.189 ;
        RECT 0.207 0.099 0.225 0.189 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.702 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.702 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.171 0.63 0.189 ;
        RECT 0.612 0.027 0.63 0.189 ;
        RECT 0.565 0.027 0.63 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.423 0.171 0.468 0.189 ;
      RECT 0.45 0.027 0.468 0.189 ;
      RECT 0.45 0.1 0.576 0.118 ;
      RECT 0.348 0.027 0.468 0.045 ;
      RECT 0.126 0.135 0.189 0.153 ;
      RECT 0.171 0.027 0.189 0.153 ;
      RECT 0.396 0.063 0.414 0.122 ;
      RECT 0.171 0.063 0.414 0.081 ;
      RECT 0.099 0.027 0.189 0.045 ;
      RECT 0.256 0.171 0.387 0.189 ;
  END
END XNOR2x2_ASAP7_6t_SL

MACRO XNOR2xp5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2xp5_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.056 0.099 0.144 0.117 ;
        RECT 0.076 0.099 0.114 0.153 ;
        RECT 0.056 0.063 0.093 0.117 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.099 0.36 0.117 ;
        RECT 0.207 0.027 0.225 0.117 ;
        RECT 0.018 0.027 0.225 0.045 ;
        RECT 0.018 0.171 0.055 0.189 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.171 0.468 0.189 ;
        RECT 0.45 0.027 0.468 0.189 ;
        RECT 0.423 0.027 0.468 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.094 0.171 0.18 0.189 ;
      RECT 0.162 0.135 0.18 0.189 ;
      RECT 0.162 0.135 0.414 0.153 ;
      RECT 0.396 0.094 0.414 0.153 ;
      RECT 0.171 0.063 0.189 0.153 ;
      RECT 0.126 0.063 0.189 0.081 ;
      RECT 0.256 0.027 0.387 0.045 ;
  END
END XNOR2xp5_ASAP7_6t_SL

MACRO XNOR2xp5f_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2xp5f_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.056 0.099 0.144 0.117 ;
        RECT 0.081 0.099 0.118 0.153 ;
        RECT 0.056 0.063 0.093 0.117 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.099 0.36 0.117 ;
        RECT 0.207 0.027 0.225 0.117 ;
        RECT 0.018 0.027 0.225 0.045 ;
        RECT 0.018 0.171 0.068 0.189 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.256 0.171 0.468 0.189 ;
        RECT 0.45 0.027 0.468 0.189 ;
        RECT 0.418 0.027 0.468 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.099 0.171 0.189 0.189 ;
      RECT 0.171 0.063 0.189 0.189 ;
      RECT 0.171 0.135 0.414 0.153 ;
      RECT 0.396 0.094 0.414 0.153 ;
      RECT 0.126 0.063 0.189 0.081 ;
      RECT 0.256 0.027 0.387 0.045 ;
  END
END XNOR2xp5f_ASAP7_6t_SL

MACRO XOR2x2_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2x2_ASAP7_6t_SL 0 0 ;
  SIZE 0.702 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.056 0.099 0.144 0.117 ;
        RECT 0.083 0.099 0.12 0.153 ;
        RECT 0.056 0.063 0.095 0.118 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.099 0.36 0.117 ;
        RECT 0.207 0.027 0.225 0.117 ;
        RECT 0.018 0.027 0.225 0.045 ;
        RECT 0.018 0.171 0.068 0.189 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.702 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.702 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.171 0.63 0.189 ;
        RECT 0.612 0.027 0.63 0.189 ;
        RECT 0.58 0.027 0.63 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.364 0.171 0.468 0.189 ;
      RECT 0.45 0.027 0.468 0.189 ;
      RECT 0.45 0.098 0.576 0.116 ;
      RECT 0.423 0.027 0.468 0.045 ;
      RECT 0.099 0.171 0.189 0.189 ;
      RECT 0.171 0.063 0.189 0.189 ;
      RECT 0.171 0.135 0.414 0.153 ;
      RECT 0.396 0.094 0.414 0.153 ;
      RECT 0.126 0.063 0.189 0.081 ;
      RECT 0.256 0.027 0.392 0.045 ;
  END
END XOR2x2_ASAP7_6t_SL

MACRO XOR2xp5_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2xp5_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.099 0.36 0.117 ;
        RECT 0.018 0.171 0.225 0.189 ;
        RECT 0.207 0.099 0.225 0.189 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.056 0.099 0.144 0.117 ;
        RECT 0.077 0.063 0.122 0.117 ;
        RECT 0.056 0.099 0.093 0.153 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.423 0.171 0.468 0.189 ;
        RECT 0.45 0.027 0.468 0.189 ;
        RECT 0.256 0.027 0.468 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.126 0.135 0.189 0.153 ;
      RECT 0.171 0.027 0.189 0.153 ;
      RECT 0.396 0.063 0.414 0.122 ;
      RECT 0.171 0.063 0.414 0.081 ;
      RECT 0.099 0.027 0.189 0.045 ;
      RECT 0.256 0.171 0.387 0.189 ;
  END
END XOR2xp5_ASAP7_6t_SL

MACRO XOR2xp5r_ASAP7_6t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2xp5r_ASAP7_6t_SL 0 0 ;
  SIZE 0.486 BY 0.216 ;
  SYMMETRY X Y ;
  SITE asap7sc6t ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.056 0.099 0.144 0.117 ;
        RECT 0.076 0.063 0.114 0.117 ;
        RECT 0.056 0.099 0.093 0.153 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.207 0.099 0.36 0.117 ;
        RECT 0.018 0.171 0.225 0.189 ;
        RECT 0.207 0.099 0.225 0.189 ;
        RECT 0.018 0.027 0.065 0.045 ;
        RECT 0.018 0.027 0.036 0.189 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.207 0.486 0.225 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 0.486 0.009 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.423 0.171 0.468 0.189 ;
        RECT 0.45 0.027 0.468 0.189 ;
        RECT 0.256 0.027 0.468 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.126 0.135 0.189 0.153 ;
      RECT 0.171 0.027 0.189 0.153 ;
      RECT 0.396 0.063 0.414 0.122 ;
      RECT 0.171 0.063 0.414 0.081 ;
      RECT 0.099 0.027 0.189 0.045 ;
      RECT 0.256 0.171 0.392 0.189 ;
  END
END XOR2xp5r_ASAP7_6t_SL

END LIBRARY
